// This is the unpowered netlist.
module Main (CLK,
    GPIO);
 input CLK;
 output [31:0] GPIO;

 wire \RAM_READ_DATA[0] ;
 wire \RAM_READ_DATA[1] ;
 wire \RAM_READ_DATA[2] ;
 wire \RAM_READ_DATA[3] ;
 wire \RAM_READ_DATA[4] ;
 wire \RAM_READ_DATA[5] ;
 wire \RAM_READ_DATA[6] ;
 wire \RAM_READ_DATA[7] ;
 wire _0000_;
 wire net254;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire net253;
 wire _0012_;
 wire clknet_leaf_0_CLK;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire net255;
 wire \cpu.ALU_OUT[0] ;
 wire \cpu.ALU_OUT[10] ;
 wire \cpu.ALU_OUT[11] ;
 wire \cpu.ALU_OUT[12] ;
 wire \cpu.ALU_OUT[13] ;
 wire \cpu.ALU_OUT[14] ;
 wire \cpu.ALU_OUT[15] ;
 wire \cpu.ALU_OUT[16] ;
 wire \cpu.ALU_OUT[17] ;
 wire \cpu.ALU_OUT[18] ;
 wire \cpu.ALU_OUT[19] ;
 wire \cpu.ALU_OUT[1] ;
 wire \cpu.ALU_OUT[20] ;
 wire \cpu.ALU_OUT[21] ;
 wire \cpu.ALU_OUT[22] ;
 wire \cpu.ALU_OUT[23] ;
 wire \cpu.ALU_OUT[24] ;
 wire \cpu.ALU_OUT[25] ;
 wire \cpu.ALU_OUT[26] ;
 wire \cpu.ALU_OUT[27] ;
 wire \cpu.ALU_OUT[28] ;
 wire \cpu.ALU_OUT[29] ;
 wire \cpu.ALU_OUT[2] ;
 wire \cpu.ALU_OUT[30] ;
 wire \cpu.ALU_OUT[31] ;
 wire \cpu.ALU_OUT[3] ;
 wire \cpu.ALU_OUT[4] ;
 wire \cpu.ALU_OUT[5] ;
 wire \cpu.ALU_OUT[6] ;
 wire \cpu.ALU_OUT[7] ;
 wire \cpu.ALU_OUT[8] ;
 wire \cpu.ALU_OUT[9] ;
 wire \cpu.ALU_OUT_MEMORY_4[0] ;
 wire \cpu.ALU_OUT_MEMORY_4[10] ;
 wire \cpu.ALU_OUT_MEMORY_4[11] ;
 wire \cpu.ALU_OUT_MEMORY_4[12] ;
 wire \cpu.ALU_OUT_MEMORY_4[13] ;
 wire \cpu.ALU_OUT_MEMORY_4[14] ;
 wire \cpu.ALU_OUT_MEMORY_4[15] ;
 wire \cpu.ALU_OUT_MEMORY_4[16] ;
 wire \cpu.ALU_OUT_MEMORY_4[17] ;
 wire \cpu.ALU_OUT_MEMORY_4[18] ;
 wire \cpu.ALU_OUT_MEMORY_4[19] ;
 wire \cpu.ALU_OUT_MEMORY_4[1] ;
 wire \cpu.ALU_OUT_MEMORY_4[20] ;
 wire \cpu.ALU_OUT_MEMORY_4[21] ;
 wire \cpu.ALU_OUT_MEMORY_4[22] ;
 wire \cpu.ALU_OUT_MEMORY_4[23] ;
 wire \cpu.ALU_OUT_MEMORY_4[24] ;
 wire \cpu.ALU_OUT_MEMORY_4[25] ;
 wire \cpu.ALU_OUT_MEMORY_4[26] ;
 wire \cpu.ALU_OUT_MEMORY_4[27] ;
 wire \cpu.ALU_OUT_MEMORY_4[28] ;
 wire \cpu.ALU_OUT_MEMORY_4[29] ;
 wire \cpu.ALU_OUT_MEMORY_4[2] ;
 wire \cpu.ALU_OUT_MEMORY_4[30] ;
 wire \cpu.ALU_OUT_MEMORY_4[31] ;
 wire \cpu.ALU_OUT_MEMORY_4[3] ;
 wire \cpu.ALU_OUT_MEMORY_4[4] ;
 wire \cpu.ALU_OUT_MEMORY_4[5] ;
 wire \cpu.ALU_OUT_MEMORY_4[6] ;
 wire \cpu.ALU_OUT_MEMORY_4[7] ;
 wire \cpu.ALU_OUT_MEMORY_4[8] ;
 wire \cpu.ALU_OUT_MEMORY_4[9] ;
 wire \cpu.INSTRUCTION_DECODE_2[0] ;
 wire \cpu.INSTRUCTION_DECODE_2[10] ;
 wire \cpu.INSTRUCTION_DECODE_2[11] ;
 wire \cpu.INSTRUCTION_DECODE_2[13] ;
 wire \cpu.INSTRUCTION_DECODE_2[16] ;
 wire \cpu.INSTRUCTION_DECODE_2[20] ;
 wire \cpu.INSTRUCTION_DECODE_2[21] ;
 wire \cpu.INSTRUCTION_DECODE_2[22] ;
 wire \cpu.INSTRUCTION_DECODE_2[4] ;
 wire \cpu.INSTRUCTION_DECODE_2[5] ;
 wire \cpu.INSTRUCTION_DECODE_2[7] ;
 wire \cpu.INSTRUCTION_DECODE_2[8] ;
 wire \cpu.INSTRUCTION_DECODE_2[9] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[0] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[10] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[11] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[13] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[16] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[20] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[21] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[22] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[4] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[5] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[7] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[8] ;
 wire \cpu.INSTRUCTION_EXECUTE_3[9] ;
 wire \cpu.INSTRUCTION_MEMORY_4[0] ;
 wire \cpu.INSTRUCTION_MEMORY_4[10] ;
 wire \cpu.INSTRUCTION_MEMORY_4[11] ;
 wire \cpu.INSTRUCTION_MEMORY_4[4] ;
 wire \cpu.INSTRUCTION_MEMORY_4[5] ;
 wire \cpu.INSTRUCTION_MEMORY_4[7] ;
 wire \cpu.INSTRUCTION_MEMORY_4[8] ;
 wire \cpu.INSTRUCTION_MEMORY_4[9] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[0] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[10] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[11] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[4] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[5] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[7] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[8] ;
 wire \cpu.INSTRUCTION_WRITEBACK_5[9] ;
 wire \cpu.PC[0] ;
 wire \cpu.PC[1] ;
 wire \cpu.PC[2] ;
 wire \cpu.PC[3] ;
 wire \cpu.PC[4] ;
 wire \cpu.PC[5] ;
 wire \cpu.PC[6] ;
 wire \cpu.PC[7] ;
 wire \cpu.PC[8] ;
 wire \cpu.PC[9] ;
 wire \cpu.PC_DECODE_2[0] ;
 wire \cpu.PC_DECODE_2[1] ;
 wire \cpu.PC_DECODE_2[2] ;
 wire \cpu.PC_DECODE_2[3] ;
 wire \cpu.PC_DECODE_2[4] ;
 wire \cpu.PC_DECODE_2[5] ;
 wire \cpu.PC_DECODE_2[6] ;
 wire \cpu.PC_DECODE_2[7] ;
 wire \cpu.PC_DECODE_2[8] ;
 wire \cpu.PC_DECODE_2[9] ;
 wire \cpu.PC_EXECUTE_3[0] ;
 wire \cpu.PC_EXECUTE_3[1] ;
 wire \cpu.PC_EXECUTE_3[2] ;
 wire \cpu.PC_EXECUTE_3[3] ;
 wire \cpu.PC_EXECUTE_3[4] ;
 wire \cpu.PC_EXECUTE_3[5] ;
 wire \cpu.PC_EXECUTE_3[6] ;
 wire \cpu.PC_EXECUTE_3[7] ;
 wire \cpu.PC_EXECUTE_3[8] ;
 wire \cpu.PC_EXECUTE_3[9] ;
 wire \cpu.PC_MEMORY_4[0] ;
 wire \cpu.PC_MEMORY_4[1] ;
 wire \cpu.PC_MEMORY_4[2] ;
 wire \cpu.PC_MEMORY_4[3] ;
 wire \cpu.PC_MEMORY_4[4] ;
 wire \cpu.PC_MEMORY_4[5] ;
 wire \cpu.PC_MEMORY_4[6] ;
 wire \cpu.PC_MEMORY_4[7] ;
 wire \cpu.PC_MEMORY_4[8] ;
 wire \cpu.PC_MEMORY_4[9] ;
 wire \cpu.R1_PIPELINE[0][1] ;
 wire \cpu.R1_PIPELINE[1][1] ;
 wire \cpu.R2_DATA[0] ;
 wire \cpu.R2_DATA[1] ;
 wire \cpu.R2_DATA[2] ;
 wire \cpu.R2_DATA[3] ;
 wire \cpu.R2_DATA[4] ;
 wire \cpu.R2_DATA[5] ;
 wire \cpu.R2_DATA[6] ;
 wire \cpu.R2_DATA[7] ;
 wire \cpu.R2_PIPELINE[0][0] ;
 wire \cpu.R2_PIPELINE[0][1] ;
 wire \cpu.R2_PIPELINE[0][2] ;
 wire \cpu.R2_PIPELINE[0][3] ;
 wire \cpu.R2_PIPELINE[1][0] ;
 wire \cpu.R2_PIPELINE[1][1] ;
 wire \cpu.R2_PIPELINE[1][2] ;
 wire \cpu.R2_PIPELINE[1][3] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[0] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[1] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[2] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[3] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[4] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[5] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[6] ;
 wire \cpu.RAM_READ_DATA_WRITEBACK_5[7] ;
 wire \cpu.RAM_WRITE_DATA[0] ;
 wire \cpu.RAM_WRITE_DATA[1] ;
 wire \cpu.RAM_WRITE_DATA[2] ;
 wire \cpu.RAM_WRITE_DATA[3] ;
 wire \cpu.RAM_WRITE_DATA[4] ;
 wire \cpu.RAM_WRITE_DATA[5] ;
 wire \cpu.RAM_WRITE_DATA[6] ;
 wire \cpu.RAM_WRITE_DATA[7] ;
 wire \cpu.RD_PIPELINE[1][0] ;
 wire \cpu.RD_PIPELINE[1][1] ;
 wire \cpu.RD_PIPELINE[1][2] ;
 wire \cpu.RD_PIPELINE[1][3] ;
 wire \cpu.RD_PIPELINE[2][0] ;
 wire \cpu.RD_PIPELINE[2][1] ;
 wire \cpu.RD_PIPELINE[2][2] ;
 wire \cpu.RD_PIPELINE[2][3] ;
 wire \cpu.RD_PIPELINE[2][4] ;
 wire \cpu.RD_PIPELINE[3][0] ;
 wire \cpu.RD_PIPELINE[3][1] ;
 wire \cpu.RD_PIPELINE[3][2] ;
 wire \cpu.RD_PIPELINE[3][3] ;
 wire \cpu.RD_PIPELINE[3][4] ;
 wire \cpu.REG_WRITE_DATA[0] ;
 wire \cpu.REG_WRITE_DATA[10] ;
 wire \cpu.REG_WRITE_DATA[11] ;
 wire \cpu.REG_WRITE_DATA[12] ;
 wire \cpu.REG_WRITE_DATA[13] ;
 wire \cpu.REG_WRITE_DATA[14] ;
 wire \cpu.REG_WRITE_DATA[15] ;
 wire \cpu.REG_WRITE_DATA[16] ;
 wire \cpu.REG_WRITE_DATA[17] ;
 wire \cpu.REG_WRITE_DATA[18] ;
 wire \cpu.REG_WRITE_DATA[19] ;
 wire \cpu.REG_WRITE_DATA[1] ;
 wire \cpu.REG_WRITE_DATA[20] ;
 wire \cpu.REG_WRITE_DATA[21] ;
 wire \cpu.REG_WRITE_DATA[22] ;
 wire \cpu.REG_WRITE_DATA[23] ;
 wire \cpu.REG_WRITE_DATA[24] ;
 wire \cpu.REG_WRITE_DATA[25] ;
 wire \cpu.REG_WRITE_DATA[26] ;
 wire \cpu.REG_WRITE_DATA[27] ;
 wire \cpu.REG_WRITE_DATA[28] ;
 wire \cpu.REG_WRITE_DATA[29] ;
 wire \cpu.REG_WRITE_DATA[2] ;
 wire \cpu.REG_WRITE_DATA[30] ;
 wire \cpu.REG_WRITE_DATA[31] ;
 wire \cpu.REG_WRITE_DATA[3] ;
 wire \cpu.REG_WRITE_DATA[4] ;
 wire \cpu.REG_WRITE_DATA[5] ;
 wire \cpu.REG_WRITE_DATA[6] ;
 wire \cpu.REG_WRITE_DATA[7] ;
 wire \cpu.REG_WRITE_DATA[8] ;
 wire \cpu.REG_WRITE_DATA[9] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[0] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[10] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[11] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[12] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[13] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[14] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[15] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[16] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[17] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[18] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[19] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[1] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[20] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[21] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[22] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[23] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[24] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[25] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[26] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[27] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[28] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[29] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[2] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[30] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[31] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[3] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[4] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[5] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[6] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[7] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[8] ;
 wire \cpu.REG_WRITE_DATA_WRITEBACK_5[9] ;
 wire \cpu.TYPE_PIPELINE[0][0] ;
 wire \cpu.TYPE_PIPELINE[0][1] ;
 wire \cpu.TYPE_PIPELINE[0][2] ;
 wire \cpu.TYPE_PIPELINE[0][3] ;
 wire \cpu.TYPE_PIPELINE[0][4] ;
 wire \cpu.TYPE_PIPELINE[1][0] ;
 wire \cpu.TYPE_PIPELINE[1][1] ;
 wire \cpu.TYPE_PIPELINE[1][2] ;
 wire \cpu.TYPE_PIPELINE[1][3] ;
 wire \cpu.TYPE_PIPELINE[1][4] ;
 wire \cpu.immediateExtractor.VALUE[0] ;
 wire \cpu.immediateExtractor.VALUE[10] ;
 wire \cpu.immediateExtractor.VALUE[11] ;
 wire \cpu.immediateExtractor.VALUE[13] ;
 wire \cpu.immediateExtractor.VALUE[16] ;
 wire \cpu.immediateExtractor.VALUE[1] ;
 wire \cpu.immediateExtractor.VALUE[20] ;
 wire \cpu.immediateExtractor.VALUE[21] ;
 wire \cpu.immediateExtractor.VALUE[22] ;
 wire \cpu.immediateExtractor.VALUE[2] ;
 wire \cpu.immediateExtractor.VALUE[31] ;
 wire \cpu.immediateExtractor.VALUE[3] ;
 wire \cpu.immediateExtractor.VALUE[4] ;
 wire \cpu.regFile.REGISTERS[0][0] ;
 wire \cpu.regFile.REGISTERS[0][10] ;
 wire \cpu.regFile.REGISTERS[0][11] ;
 wire \cpu.regFile.REGISTERS[0][12] ;
 wire \cpu.regFile.REGISTERS[0][13] ;
 wire \cpu.regFile.REGISTERS[0][14] ;
 wire \cpu.regFile.REGISTERS[0][15] ;
 wire \cpu.regFile.REGISTERS[0][16] ;
 wire \cpu.regFile.REGISTERS[0][17] ;
 wire \cpu.regFile.REGISTERS[0][18] ;
 wire \cpu.regFile.REGISTERS[0][19] ;
 wire \cpu.regFile.REGISTERS[0][1] ;
 wire \cpu.regFile.REGISTERS[0][20] ;
 wire \cpu.regFile.REGISTERS[0][21] ;
 wire \cpu.regFile.REGISTERS[0][22] ;
 wire \cpu.regFile.REGISTERS[0][23] ;
 wire \cpu.regFile.REGISTERS[0][24] ;
 wire \cpu.regFile.REGISTERS[0][25] ;
 wire \cpu.regFile.REGISTERS[0][26] ;
 wire \cpu.regFile.REGISTERS[0][27] ;
 wire \cpu.regFile.REGISTERS[0][28] ;
 wire \cpu.regFile.REGISTERS[0][29] ;
 wire \cpu.regFile.REGISTERS[0][2] ;
 wire \cpu.regFile.REGISTERS[0][30] ;
 wire \cpu.regFile.REGISTERS[0][31] ;
 wire \cpu.regFile.REGISTERS[0][3] ;
 wire \cpu.regFile.REGISTERS[0][4] ;
 wire \cpu.regFile.REGISTERS[0][5] ;
 wire \cpu.regFile.REGISTERS[0][6] ;
 wire \cpu.regFile.REGISTERS[0][7] ;
 wire \cpu.regFile.REGISTERS[0][8] ;
 wire \cpu.regFile.REGISTERS[0][9] ;
 wire \cpu.regFile.REGISTERS[10][0] ;
 wire \cpu.regFile.REGISTERS[10][10] ;
 wire \cpu.regFile.REGISTERS[10][11] ;
 wire \cpu.regFile.REGISTERS[10][12] ;
 wire \cpu.regFile.REGISTERS[10][13] ;
 wire \cpu.regFile.REGISTERS[10][14] ;
 wire \cpu.regFile.REGISTERS[10][15] ;
 wire \cpu.regFile.REGISTERS[10][16] ;
 wire \cpu.regFile.REGISTERS[10][17] ;
 wire \cpu.regFile.REGISTERS[10][18] ;
 wire \cpu.regFile.REGISTERS[10][19] ;
 wire \cpu.regFile.REGISTERS[10][1] ;
 wire \cpu.regFile.REGISTERS[10][20] ;
 wire \cpu.regFile.REGISTERS[10][21] ;
 wire \cpu.regFile.REGISTERS[10][22] ;
 wire \cpu.regFile.REGISTERS[10][23] ;
 wire \cpu.regFile.REGISTERS[10][24] ;
 wire \cpu.regFile.REGISTERS[10][25] ;
 wire \cpu.regFile.REGISTERS[10][26] ;
 wire \cpu.regFile.REGISTERS[10][27] ;
 wire \cpu.regFile.REGISTERS[10][28] ;
 wire \cpu.regFile.REGISTERS[10][29] ;
 wire \cpu.regFile.REGISTERS[10][2] ;
 wire \cpu.regFile.REGISTERS[10][30] ;
 wire \cpu.regFile.REGISTERS[10][31] ;
 wire \cpu.regFile.REGISTERS[10][3] ;
 wire \cpu.regFile.REGISTERS[10][4] ;
 wire \cpu.regFile.REGISTERS[10][5] ;
 wire \cpu.regFile.REGISTERS[10][6] ;
 wire \cpu.regFile.REGISTERS[10][7] ;
 wire \cpu.regFile.REGISTERS[10][8] ;
 wire \cpu.regFile.REGISTERS[10][9] ;
 wire \cpu.regFile.REGISTERS[11][0] ;
 wire \cpu.regFile.REGISTERS[11][10] ;
 wire \cpu.regFile.REGISTERS[11][11] ;
 wire \cpu.regFile.REGISTERS[11][12] ;
 wire \cpu.regFile.REGISTERS[11][13] ;
 wire \cpu.regFile.REGISTERS[11][14] ;
 wire \cpu.regFile.REGISTERS[11][15] ;
 wire \cpu.regFile.REGISTERS[11][16] ;
 wire \cpu.regFile.REGISTERS[11][17] ;
 wire \cpu.regFile.REGISTERS[11][18] ;
 wire \cpu.regFile.REGISTERS[11][19] ;
 wire \cpu.regFile.REGISTERS[11][1] ;
 wire \cpu.regFile.REGISTERS[11][20] ;
 wire \cpu.regFile.REGISTERS[11][21] ;
 wire \cpu.regFile.REGISTERS[11][22] ;
 wire \cpu.regFile.REGISTERS[11][23] ;
 wire \cpu.regFile.REGISTERS[11][24] ;
 wire \cpu.regFile.REGISTERS[11][25] ;
 wire \cpu.regFile.REGISTERS[11][26] ;
 wire \cpu.regFile.REGISTERS[11][27] ;
 wire \cpu.regFile.REGISTERS[11][28] ;
 wire \cpu.regFile.REGISTERS[11][29] ;
 wire \cpu.regFile.REGISTERS[11][2] ;
 wire \cpu.regFile.REGISTERS[11][30] ;
 wire \cpu.regFile.REGISTERS[11][31] ;
 wire \cpu.regFile.REGISTERS[11][3] ;
 wire \cpu.regFile.REGISTERS[11][4] ;
 wire \cpu.regFile.REGISTERS[11][5] ;
 wire \cpu.regFile.REGISTERS[11][6] ;
 wire \cpu.regFile.REGISTERS[11][7] ;
 wire \cpu.regFile.REGISTERS[11][8] ;
 wire \cpu.regFile.REGISTERS[11][9] ;
 wire \cpu.regFile.REGISTERS[12][0] ;
 wire \cpu.regFile.REGISTERS[12][10] ;
 wire \cpu.regFile.REGISTERS[12][11] ;
 wire \cpu.regFile.REGISTERS[12][12] ;
 wire \cpu.regFile.REGISTERS[12][13] ;
 wire \cpu.regFile.REGISTERS[12][14] ;
 wire \cpu.regFile.REGISTERS[12][15] ;
 wire \cpu.regFile.REGISTERS[12][16] ;
 wire \cpu.regFile.REGISTERS[12][17] ;
 wire \cpu.regFile.REGISTERS[12][18] ;
 wire \cpu.regFile.REGISTERS[12][19] ;
 wire \cpu.regFile.REGISTERS[12][1] ;
 wire \cpu.regFile.REGISTERS[12][20] ;
 wire \cpu.regFile.REGISTERS[12][21] ;
 wire \cpu.regFile.REGISTERS[12][22] ;
 wire \cpu.regFile.REGISTERS[12][23] ;
 wire \cpu.regFile.REGISTERS[12][24] ;
 wire \cpu.regFile.REGISTERS[12][25] ;
 wire \cpu.regFile.REGISTERS[12][26] ;
 wire \cpu.regFile.REGISTERS[12][27] ;
 wire \cpu.regFile.REGISTERS[12][28] ;
 wire \cpu.regFile.REGISTERS[12][29] ;
 wire \cpu.regFile.REGISTERS[12][2] ;
 wire \cpu.regFile.REGISTERS[12][30] ;
 wire \cpu.regFile.REGISTERS[12][31] ;
 wire \cpu.regFile.REGISTERS[12][3] ;
 wire \cpu.regFile.REGISTERS[12][4] ;
 wire \cpu.regFile.REGISTERS[12][5] ;
 wire \cpu.regFile.REGISTERS[12][6] ;
 wire \cpu.regFile.REGISTERS[12][7] ;
 wire \cpu.regFile.REGISTERS[12][8] ;
 wire \cpu.regFile.REGISTERS[12][9] ;
 wire \cpu.regFile.REGISTERS[13][0] ;
 wire \cpu.regFile.REGISTERS[13][10] ;
 wire \cpu.regFile.REGISTERS[13][11] ;
 wire \cpu.regFile.REGISTERS[13][12] ;
 wire \cpu.regFile.REGISTERS[13][13] ;
 wire \cpu.regFile.REGISTERS[13][14] ;
 wire \cpu.regFile.REGISTERS[13][15] ;
 wire \cpu.regFile.REGISTERS[13][16] ;
 wire \cpu.regFile.REGISTERS[13][17] ;
 wire \cpu.regFile.REGISTERS[13][18] ;
 wire \cpu.regFile.REGISTERS[13][19] ;
 wire \cpu.regFile.REGISTERS[13][1] ;
 wire \cpu.regFile.REGISTERS[13][20] ;
 wire \cpu.regFile.REGISTERS[13][21] ;
 wire \cpu.regFile.REGISTERS[13][22] ;
 wire \cpu.regFile.REGISTERS[13][23] ;
 wire \cpu.regFile.REGISTERS[13][24] ;
 wire \cpu.regFile.REGISTERS[13][25] ;
 wire \cpu.regFile.REGISTERS[13][26] ;
 wire \cpu.regFile.REGISTERS[13][27] ;
 wire \cpu.regFile.REGISTERS[13][28] ;
 wire \cpu.regFile.REGISTERS[13][29] ;
 wire \cpu.regFile.REGISTERS[13][2] ;
 wire \cpu.regFile.REGISTERS[13][30] ;
 wire \cpu.regFile.REGISTERS[13][31] ;
 wire \cpu.regFile.REGISTERS[13][3] ;
 wire \cpu.regFile.REGISTERS[13][4] ;
 wire \cpu.regFile.REGISTERS[13][5] ;
 wire \cpu.regFile.REGISTERS[13][6] ;
 wire \cpu.regFile.REGISTERS[13][7] ;
 wire \cpu.regFile.REGISTERS[13][8] ;
 wire \cpu.regFile.REGISTERS[13][9] ;
 wire \cpu.regFile.REGISTERS[14][0] ;
 wire \cpu.regFile.REGISTERS[14][10] ;
 wire \cpu.regFile.REGISTERS[14][11] ;
 wire \cpu.regFile.REGISTERS[14][12] ;
 wire \cpu.regFile.REGISTERS[14][13] ;
 wire \cpu.regFile.REGISTERS[14][14] ;
 wire \cpu.regFile.REGISTERS[14][15] ;
 wire \cpu.regFile.REGISTERS[14][16] ;
 wire \cpu.regFile.REGISTERS[14][17] ;
 wire \cpu.regFile.REGISTERS[14][18] ;
 wire \cpu.regFile.REGISTERS[14][19] ;
 wire \cpu.regFile.REGISTERS[14][1] ;
 wire \cpu.regFile.REGISTERS[14][20] ;
 wire \cpu.regFile.REGISTERS[14][21] ;
 wire \cpu.regFile.REGISTERS[14][22] ;
 wire \cpu.regFile.REGISTERS[14][23] ;
 wire \cpu.regFile.REGISTERS[14][24] ;
 wire \cpu.regFile.REGISTERS[14][25] ;
 wire \cpu.regFile.REGISTERS[14][26] ;
 wire \cpu.regFile.REGISTERS[14][27] ;
 wire \cpu.regFile.REGISTERS[14][28] ;
 wire \cpu.regFile.REGISTERS[14][29] ;
 wire \cpu.regFile.REGISTERS[14][2] ;
 wire \cpu.regFile.REGISTERS[14][30] ;
 wire \cpu.regFile.REGISTERS[14][31] ;
 wire \cpu.regFile.REGISTERS[14][3] ;
 wire \cpu.regFile.REGISTERS[14][4] ;
 wire \cpu.regFile.REGISTERS[14][5] ;
 wire \cpu.regFile.REGISTERS[14][6] ;
 wire \cpu.regFile.REGISTERS[14][7] ;
 wire \cpu.regFile.REGISTERS[14][8] ;
 wire \cpu.regFile.REGISTERS[14][9] ;
 wire \cpu.regFile.REGISTERS[15][0] ;
 wire \cpu.regFile.REGISTERS[15][10] ;
 wire \cpu.regFile.REGISTERS[15][11] ;
 wire \cpu.regFile.REGISTERS[15][12] ;
 wire \cpu.regFile.REGISTERS[15][13] ;
 wire \cpu.regFile.REGISTERS[15][14] ;
 wire \cpu.regFile.REGISTERS[15][15] ;
 wire \cpu.regFile.REGISTERS[15][16] ;
 wire \cpu.regFile.REGISTERS[15][17] ;
 wire \cpu.regFile.REGISTERS[15][18] ;
 wire \cpu.regFile.REGISTERS[15][19] ;
 wire \cpu.regFile.REGISTERS[15][1] ;
 wire \cpu.regFile.REGISTERS[15][20] ;
 wire \cpu.regFile.REGISTERS[15][21] ;
 wire \cpu.regFile.REGISTERS[15][22] ;
 wire \cpu.regFile.REGISTERS[15][23] ;
 wire \cpu.regFile.REGISTERS[15][24] ;
 wire \cpu.regFile.REGISTERS[15][25] ;
 wire \cpu.regFile.REGISTERS[15][26] ;
 wire \cpu.regFile.REGISTERS[15][27] ;
 wire \cpu.regFile.REGISTERS[15][28] ;
 wire \cpu.regFile.REGISTERS[15][29] ;
 wire \cpu.regFile.REGISTERS[15][2] ;
 wire \cpu.regFile.REGISTERS[15][30] ;
 wire \cpu.regFile.REGISTERS[15][31] ;
 wire \cpu.regFile.REGISTERS[15][3] ;
 wire \cpu.regFile.REGISTERS[15][4] ;
 wire \cpu.regFile.REGISTERS[15][5] ;
 wire \cpu.regFile.REGISTERS[15][6] ;
 wire \cpu.regFile.REGISTERS[15][7] ;
 wire \cpu.regFile.REGISTERS[15][8] ;
 wire \cpu.regFile.REGISTERS[15][9] ;
 wire \cpu.regFile.REGISTERS[1][0] ;
 wire \cpu.regFile.REGISTERS[1][10] ;
 wire \cpu.regFile.REGISTERS[1][11] ;
 wire \cpu.regFile.REGISTERS[1][12] ;
 wire \cpu.regFile.REGISTERS[1][13] ;
 wire \cpu.regFile.REGISTERS[1][14] ;
 wire \cpu.regFile.REGISTERS[1][15] ;
 wire \cpu.regFile.REGISTERS[1][16] ;
 wire \cpu.regFile.REGISTERS[1][17] ;
 wire \cpu.regFile.REGISTERS[1][18] ;
 wire \cpu.regFile.REGISTERS[1][19] ;
 wire \cpu.regFile.REGISTERS[1][1] ;
 wire \cpu.regFile.REGISTERS[1][20] ;
 wire \cpu.regFile.REGISTERS[1][21] ;
 wire \cpu.regFile.REGISTERS[1][22] ;
 wire \cpu.regFile.REGISTERS[1][23] ;
 wire \cpu.regFile.REGISTERS[1][24] ;
 wire \cpu.regFile.REGISTERS[1][25] ;
 wire \cpu.regFile.REGISTERS[1][26] ;
 wire \cpu.regFile.REGISTERS[1][27] ;
 wire \cpu.regFile.REGISTERS[1][28] ;
 wire \cpu.regFile.REGISTERS[1][29] ;
 wire \cpu.regFile.REGISTERS[1][2] ;
 wire \cpu.regFile.REGISTERS[1][30] ;
 wire \cpu.regFile.REGISTERS[1][31] ;
 wire \cpu.regFile.REGISTERS[1][3] ;
 wire \cpu.regFile.REGISTERS[1][4] ;
 wire \cpu.regFile.REGISTERS[1][5] ;
 wire \cpu.regFile.REGISTERS[1][6] ;
 wire \cpu.regFile.REGISTERS[1][7] ;
 wire \cpu.regFile.REGISTERS[1][8] ;
 wire \cpu.regFile.REGISTERS[1][9] ;
 wire \cpu.regFile.REGISTERS[2][0] ;
 wire \cpu.regFile.REGISTERS[2][10] ;
 wire \cpu.regFile.REGISTERS[2][11] ;
 wire \cpu.regFile.REGISTERS[2][12] ;
 wire \cpu.regFile.REGISTERS[2][13] ;
 wire \cpu.regFile.REGISTERS[2][14] ;
 wire \cpu.regFile.REGISTERS[2][15] ;
 wire \cpu.regFile.REGISTERS[2][16] ;
 wire \cpu.regFile.REGISTERS[2][17] ;
 wire \cpu.regFile.REGISTERS[2][18] ;
 wire \cpu.regFile.REGISTERS[2][19] ;
 wire \cpu.regFile.REGISTERS[2][1] ;
 wire \cpu.regFile.REGISTERS[2][20] ;
 wire \cpu.regFile.REGISTERS[2][21] ;
 wire \cpu.regFile.REGISTERS[2][22] ;
 wire \cpu.regFile.REGISTERS[2][23] ;
 wire \cpu.regFile.REGISTERS[2][24] ;
 wire \cpu.regFile.REGISTERS[2][25] ;
 wire \cpu.regFile.REGISTERS[2][26] ;
 wire \cpu.regFile.REGISTERS[2][27] ;
 wire \cpu.regFile.REGISTERS[2][28] ;
 wire \cpu.regFile.REGISTERS[2][29] ;
 wire \cpu.regFile.REGISTERS[2][2] ;
 wire \cpu.regFile.REGISTERS[2][30] ;
 wire \cpu.regFile.REGISTERS[2][31] ;
 wire \cpu.regFile.REGISTERS[2][3] ;
 wire \cpu.regFile.REGISTERS[2][4] ;
 wire \cpu.regFile.REGISTERS[2][5] ;
 wire \cpu.regFile.REGISTERS[2][6] ;
 wire \cpu.regFile.REGISTERS[2][7] ;
 wire \cpu.regFile.REGISTERS[2][8] ;
 wire \cpu.regFile.REGISTERS[2][9] ;
 wire \cpu.regFile.REGISTERS[3][0] ;
 wire \cpu.regFile.REGISTERS[3][10] ;
 wire \cpu.regFile.REGISTERS[3][11] ;
 wire \cpu.regFile.REGISTERS[3][12] ;
 wire \cpu.regFile.REGISTERS[3][13] ;
 wire \cpu.regFile.REGISTERS[3][14] ;
 wire \cpu.regFile.REGISTERS[3][15] ;
 wire \cpu.regFile.REGISTERS[3][16] ;
 wire \cpu.regFile.REGISTERS[3][17] ;
 wire \cpu.regFile.REGISTERS[3][18] ;
 wire \cpu.regFile.REGISTERS[3][19] ;
 wire \cpu.regFile.REGISTERS[3][1] ;
 wire \cpu.regFile.REGISTERS[3][20] ;
 wire \cpu.regFile.REGISTERS[3][21] ;
 wire \cpu.regFile.REGISTERS[3][22] ;
 wire \cpu.regFile.REGISTERS[3][23] ;
 wire \cpu.regFile.REGISTERS[3][24] ;
 wire \cpu.regFile.REGISTERS[3][25] ;
 wire \cpu.regFile.REGISTERS[3][26] ;
 wire \cpu.regFile.REGISTERS[3][27] ;
 wire \cpu.regFile.REGISTERS[3][28] ;
 wire \cpu.regFile.REGISTERS[3][29] ;
 wire \cpu.regFile.REGISTERS[3][2] ;
 wire \cpu.regFile.REGISTERS[3][30] ;
 wire \cpu.regFile.REGISTERS[3][31] ;
 wire \cpu.regFile.REGISTERS[3][3] ;
 wire \cpu.regFile.REGISTERS[3][4] ;
 wire \cpu.regFile.REGISTERS[3][5] ;
 wire \cpu.regFile.REGISTERS[3][6] ;
 wire \cpu.regFile.REGISTERS[3][7] ;
 wire \cpu.regFile.REGISTERS[3][8] ;
 wire \cpu.regFile.REGISTERS[3][9] ;
 wire \cpu.regFile.REGISTERS[4][0] ;
 wire \cpu.regFile.REGISTERS[4][10] ;
 wire \cpu.regFile.REGISTERS[4][11] ;
 wire \cpu.regFile.REGISTERS[4][12] ;
 wire \cpu.regFile.REGISTERS[4][13] ;
 wire \cpu.regFile.REGISTERS[4][14] ;
 wire \cpu.regFile.REGISTERS[4][15] ;
 wire \cpu.regFile.REGISTERS[4][16] ;
 wire \cpu.regFile.REGISTERS[4][17] ;
 wire \cpu.regFile.REGISTERS[4][18] ;
 wire \cpu.regFile.REGISTERS[4][19] ;
 wire \cpu.regFile.REGISTERS[4][1] ;
 wire \cpu.regFile.REGISTERS[4][20] ;
 wire \cpu.regFile.REGISTERS[4][21] ;
 wire \cpu.regFile.REGISTERS[4][22] ;
 wire \cpu.regFile.REGISTERS[4][23] ;
 wire \cpu.regFile.REGISTERS[4][24] ;
 wire \cpu.regFile.REGISTERS[4][25] ;
 wire \cpu.regFile.REGISTERS[4][26] ;
 wire \cpu.regFile.REGISTERS[4][27] ;
 wire \cpu.regFile.REGISTERS[4][28] ;
 wire \cpu.regFile.REGISTERS[4][29] ;
 wire \cpu.regFile.REGISTERS[4][2] ;
 wire \cpu.regFile.REGISTERS[4][30] ;
 wire \cpu.regFile.REGISTERS[4][31] ;
 wire \cpu.regFile.REGISTERS[4][3] ;
 wire \cpu.regFile.REGISTERS[4][4] ;
 wire \cpu.regFile.REGISTERS[4][5] ;
 wire \cpu.regFile.REGISTERS[4][6] ;
 wire \cpu.regFile.REGISTERS[4][7] ;
 wire \cpu.regFile.REGISTERS[4][8] ;
 wire \cpu.regFile.REGISTERS[4][9] ;
 wire \cpu.regFile.REGISTERS[5][0] ;
 wire \cpu.regFile.REGISTERS[5][10] ;
 wire \cpu.regFile.REGISTERS[5][11] ;
 wire \cpu.regFile.REGISTERS[5][12] ;
 wire \cpu.regFile.REGISTERS[5][13] ;
 wire \cpu.regFile.REGISTERS[5][14] ;
 wire \cpu.regFile.REGISTERS[5][15] ;
 wire \cpu.regFile.REGISTERS[5][16] ;
 wire \cpu.regFile.REGISTERS[5][17] ;
 wire \cpu.regFile.REGISTERS[5][18] ;
 wire \cpu.regFile.REGISTERS[5][19] ;
 wire \cpu.regFile.REGISTERS[5][1] ;
 wire \cpu.regFile.REGISTERS[5][20] ;
 wire \cpu.regFile.REGISTERS[5][21] ;
 wire \cpu.regFile.REGISTERS[5][22] ;
 wire \cpu.regFile.REGISTERS[5][23] ;
 wire \cpu.regFile.REGISTERS[5][24] ;
 wire \cpu.regFile.REGISTERS[5][25] ;
 wire \cpu.regFile.REGISTERS[5][26] ;
 wire \cpu.regFile.REGISTERS[5][27] ;
 wire \cpu.regFile.REGISTERS[5][28] ;
 wire \cpu.regFile.REGISTERS[5][29] ;
 wire \cpu.regFile.REGISTERS[5][2] ;
 wire \cpu.regFile.REGISTERS[5][30] ;
 wire \cpu.regFile.REGISTERS[5][31] ;
 wire \cpu.regFile.REGISTERS[5][3] ;
 wire \cpu.regFile.REGISTERS[5][4] ;
 wire \cpu.regFile.REGISTERS[5][5] ;
 wire \cpu.regFile.REGISTERS[5][6] ;
 wire \cpu.regFile.REGISTERS[5][7] ;
 wire \cpu.regFile.REGISTERS[5][8] ;
 wire \cpu.regFile.REGISTERS[5][9] ;
 wire \cpu.regFile.REGISTERS[6][0] ;
 wire \cpu.regFile.REGISTERS[6][10] ;
 wire \cpu.regFile.REGISTERS[6][11] ;
 wire \cpu.regFile.REGISTERS[6][12] ;
 wire \cpu.regFile.REGISTERS[6][13] ;
 wire \cpu.regFile.REGISTERS[6][14] ;
 wire \cpu.regFile.REGISTERS[6][15] ;
 wire \cpu.regFile.REGISTERS[6][16] ;
 wire \cpu.regFile.REGISTERS[6][17] ;
 wire \cpu.regFile.REGISTERS[6][18] ;
 wire \cpu.regFile.REGISTERS[6][19] ;
 wire \cpu.regFile.REGISTERS[6][1] ;
 wire \cpu.regFile.REGISTERS[6][20] ;
 wire \cpu.regFile.REGISTERS[6][21] ;
 wire \cpu.regFile.REGISTERS[6][22] ;
 wire \cpu.regFile.REGISTERS[6][23] ;
 wire \cpu.regFile.REGISTERS[6][24] ;
 wire \cpu.regFile.REGISTERS[6][25] ;
 wire \cpu.regFile.REGISTERS[6][26] ;
 wire \cpu.regFile.REGISTERS[6][27] ;
 wire \cpu.regFile.REGISTERS[6][28] ;
 wire \cpu.regFile.REGISTERS[6][29] ;
 wire \cpu.regFile.REGISTERS[6][2] ;
 wire \cpu.regFile.REGISTERS[6][30] ;
 wire \cpu.regFile.REGISTERS[6][31] ;
 wire \cpu.regFile.REGISTERS[6][3] ;
 wire \cpu.regFile.REGISTERS[6][4] ;
 wire \cpu.regFile.REGISTERS[6][5] ;
 wire \cpu.regFile.REGISTERS[6][6] ;
 wire \cpu.regFile.REGISTERS[6][7] ;
 wire \cpu.regFile.REGISTERS[6][8] ;
 wire \cpu.regFile.REGISTERS[6][9] ;
 wire \cpu.regFile.REGISTERS[7][0] ;
 wire \cpu.regFile.REGISTERS[7][10] ;
 wire \cpu.regFile.REGISTERS[7][11] ;
 wire \cpu.regFile.REGISTERS[7][12] ;
 wire \cpu.regFile.REGISTERS[7][13] ;
 wire \cpu.regFile.REGISTERS[7][14] ;
 wire \cpu.regFile.REGISTERS[7][15] ;
 wire \cpu.regFile.REGISTERS[7][16] ;
 wire \cpu.regFile.REGISTERS[7][17] ;
 wire \cpu.regFile.REGISTERS[7][18] ;
 wire \cpu.regFile.REGISTERS[7][19] ;
 wire \cpu.regFile.REGISTERS[7][1] ;
 wire \cpu.regFile.REGISTERS[7][20] ;
 wire \cpu.regFile.REGISTERS[7][21] ;
 wire \cpu.regFile.REGISTERS[7][22] ;
 wire \cpu.regFile.REGISTERS[7][23] ;
 wire \cpu.regFile.REGISTERS[7][24] ;
 wire \cpu.regFile.REGISTERS[7][25] ;
 wire \cpu.regFile.REGISTERS[7][26] ;
 wire \cpu.regFile.REGISTERS[7][27] ;
 wire \cpu.regFile.REGISTERS[7][28] ;
 wire \cpu.regFile.REGISTERS[7][29] ;
 wire \cpu.regFile.REGISTERS[7][2] ;
 wire \cpu.regFile.REGISTERS[7][30] ;
 wire \cpu.regFile.REGISTERS[7][31] ;
 wire \cpu.regFile.REGISTERS[7][3] ;
 wire \cpu.regFile.REGISTERS[7][4] ;
 wire \cpu.regFile.REGISTERS[7][5] ;
 wire \cpu.regFile.REGISTERS[7][6] ;
 wire \cpu.regFile.REGISTERS[7][7] ;
 wire \cpu.regFile.REGISTERS[7][8] ;
 wire \cpu.regFile.REGISTERS[7][9] ;
 wire \cpu.regFile.REGISTERS[8][0] ;
 wire \cpu.regFile.REGISTERS[8][10] ;
 wire \cpu.regFile.REGISTERS[8][11] ;
 wire \cpu.regFile.REGISTERS[8][12] ;
 wire \cpu.regFile.REGISTERS[8][13] ;
 wire \cpu.regFile.REGISTERS[8][14] ;
 wire \cpu.regFile.REGISTERS[8][15] ;
 wire \cpu.regFile.REGISTERS[8][16] ;
 wire \cpu.regFile.REGISTERS[8][17] ;
 wire \cpu.regFile.REGISTERS[8][18] ;
 wire \cpu.regFile.REGISTERS[8][19] ;
 wire \cpu.regFile.REGISTERS[8][1] ;
 wire \cpu.regFile.REGISTERS[8][20] ;
 wire \cpu.regFile.REGISTERS[8][21] ;
 wire \cpu.regFile.REGISTERS[8][22] ;
 wire \cpu.regFile.REGISTERS[8][23] ;
 wire \cpu.regFile.REGISTERS[8][24] ;
 wire \cpu.regFile.REGISTERS[8][25] ;
 wire \cpu.regFile.REGISTERS[8][26] ;
 wire \cpu.regFile.REGISTERS[8][27] ;
 wire \cpu.regFile.REGISTERS[8][28] ;
 wire \cpu.regFile.REGISTERS[8][29] ;
 wire \cpu.regFile.REGISTERS[8][2] ;
 wire \cpu.regFile.REGISTERS[8][30] ;
 wire \cpu.regFile.REGISTERS[8][31] ;
 wire \cpu.regFile.REGISTERS[8][3] ;
 wire \cpu.regFile.REGISTERS[8][4] ;
 wire \cpu.regFile.REGISTERS[8][5] ;
 wire \cpu.regFile.REGISTERS[8][6] ;
 wire \cpu.regFile.REGISTERS[8][7] ;
 wire \cpu.regFile.REGISTERS[8][8] ;
 wire \cpu.regFile.REGISTERS[8][9] ;
 wire \cpu.regFile.REGISTERS[9][0] ;
 wire \cpu.regFile.REGISTERS[9][10] ;
 wire \cpu.regFile.REGISTERS[9][11] ;
 wire \cpu.regFile.REGISTERS[9][12] ;
 wire \cpu.regFile.REGISTERS[9][13] ;
 wire \cpu.regFile.REGISTERS[9][14] ;
 wire \cpu.regFile.REGISTERS[9][15] ;
 wire \cpu.regFile.REGISTERS[9][16] ;
 wire \cpu.regFile.REGISTERS[9][17] ;
 wire \cpu.regFile.REGISTERS[9][18] ;
 wire \cpu.regFile.REGISTERS[9][19] ;
 wire \cpu.regFile.REGISTERS[9][1] ;
 wire \cpu.regFile.REGISTERS[9][20] ;
 wire \cpu.regFile.REGISTERS[9][21] ;
 wire \cpu.regFile.REGISTERS[9][22] ;
 wire \cpu.regFile.REGISTERS[9][23] ;
 wire \cpu.regFile.REGISTERS[9][24] ;
 wire \cpu.regFile.REGISTERS[9][25] ;
 wire \cpu.regFile.REGISTERS[9][26] ;
 wire \cpu.regFile.REGISTERS[9][27] ;
 wire \cpu.regFile.REGISTERS[9][28] ;
 wire \cpu.regFile.REGISTERS[9][29] ;
 wire \cpu.regFile.REGISTERS[9][2] ;
 wire \cpu.regFile.REGISTERS[9][30] ;
 wire \cpu.regFile.REGISTERS[9][31] ;
 wire \cpu.regFile.REGISTERS[9][3] ;
 wire \cpu.regFile.REGISTERS[9][4] ;
 wire \cpu.regFile.REGISTERS[9][5] ;
 wire \cpu.regFile.REGISTERS[9][6] ;
 wire \cpu.regFile.REGISTERS[9][7] ;
 wire \cpu.regFile.REGISTERS[9][8] ;
 wire \cpu.regFile.REGISTERS[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire clknet_leaf_1_CLK;
 wire clknet_leaf_2_CLK;
 wire clknet_leaf_3_CLK;
 wire clknet_leaf_4_CLK;
 wire clknet_leaf_5_CLK;
 wire clknet_leaf_7_CLK;
 wire clknet_leaf_8_CLK;
 wire clknet_leaf_9_CLK;
 wire clknet_leaf_10_CLK;
 wire clknet_leaf_11_CLK;
 wire clknet_leaf_12_CLK;
 wire clknet_leaf_13_CLK;
 wire clknet_leaf_14_CLK;
 wire clknet_leaf_15_CLK;
 wire clknet_leaf_16_CLK;
 wire clknet_leaf_17_CLK;
 wire clknet_leaf_18_CLK;
 wire clknet_leaf_19_CLK;
 wire clknet_leaf_21_CLK;
 wire clknet_leaf_23_CLK;
 wire clknet_leaf_24_CLK;
 wire clknet_leaf_25_CLK;
 wire clknet_leaf_26_CLK;
 wire clknet_leaf_28_CLK;
 wire clknet_leaf_29_CLK;
 wire clknet_leaf_30_CLK;
 wire clknet_leaf_31_CLK;
 wire clknet_leaf_32_CLK;
 wire clknet_leaf_33_CLK;
 wire clknet_leaf_34_CLK;
 wire clknet_leaf_35_CLK;
 wire clknet_leaf_36_CLK;
 wire clknet_leaf_37_CLK;
 wire clknet_leaf_38_CLK;
 wire clknet_leaf_39_CLK;
 wire clknet_leaf_40_CLK;
 wire clknet_leaf_41_CLK;
 wire clknet_leaf_42_CLK;
 wire clknet_leaf_43_CLK;
 wire clknet_0_CLK;
 wire clknet_2_0__leaf_CLK;
 wire clknet_2_1__leaf_CLK;
 wire clknet_2_2__leaf_CLK;
 wire clknet_2_3__leaf_CLK;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;

 sky130_fd_sc_hd__buf_4 _1662_ (.A(\cpu.INSTRUCTION_EXECUTE_3[11] ),
    .X(_0207_));
 sky130_fd_sc_hd__and3b_1 _1663_ (.A_N(\cpu.INSTRUCTION_EXECUTE_3[4] ),
    .B(\cpu.INSTRUCTION_EXECUTE_3[5] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[0] ),
    .X(_0208_));
 sky130_fd_sc_hd__buf_2 _1664_ (.A(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1665_ (.A(_0207_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__buf_4 _1666_ (.A(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__clkinv_2 _1667_ (.A(_0211_),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _1668_ (.A(\cpu.INSTRUCTION_DECODE_2[4] ),
    .Y(_0212_));
 sky130_fd_sc_hd__and4_1 _1669_ (.A(\cpu.INSTRUCTION_DECODE_2[0] ),
    .B(_0212_),
    .C(\cpu.INSTRUCTION_DECODE_2[5] ),
    .D(\cpu.INSTRUCTION_DECODE_2[11] ),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _1670_ (.A(_0206_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__buf_2 _1671_ (.A(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__and2b_1 _1672_ (.A_N(\cpu.PC[3] ),
    .B(\cpu.PC[2] ),
    .X(_0216_));
 sky130_fd_sc_hd__and2b_1 _1673_ (.A_N(\cpu.PC[2] ),
    .B(\cpu.PC[3] ),
    .X(_0217_));
 sky130_fd_sc_hd__or3b_1 _1674_ (.A(\cpu.PC[5] ),
    .B(_0217_),
    .C_N(\cpu.PC[4] ),
    .X(_0218_));
 sky130_fd_sc_hd__or2_1 _1675_ (.A(_0216_),
    .B(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_0215_),
    .B(_0219_),
    .Y(_0002_));
 sky130_fd_sc_hd__or4b_1 _1677_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[5] ),
    .B(\cpu.INSTRUCTION_WRITEBACK_5[4] ),
    .C(\cpu.INSTRUCTION_WRITEBACK_5[11] ),
    .D_N(\cpu.INSTRUCTION_WRITEBACK_5[0] ),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_4 _1678_ (.A(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[1] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[1] ),
    .S(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _1680_ (.A(_0222_),
    .X(\cpu.REG_WRITE_DATA[1] ));
 sky130_fd_sc_hd__or4_1 _1681_ (.A(\cpu.TYPE_PIPELINE[1][3] ),
    .B(\cpu.TYPE_PIPELINE[1][1] ),
    .C(\cpu.TYPE_PIPELINE[1][2] ),
    .D(\cpu.TYPE_PIPELINE[1][4] ),
    .X(_0223_));
 sky130_fd_sc_hd__or4_1 _1682_ (.A(\cpu.R2_PIPELINE[1][3] ),
    .B(\cpu.R2_PIPELINE[1][1] ),
    .C(\cpu.R2_PIPELINE[1][0] ),
    .D(\cpu.R2_PIPELINE[1][2] ),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_2 _1683_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _1684_ (.A(\cpu.R2_PIPELINE[1][0] ),
    .Y(_0226_));
 sky130_fd_sc_hd__or2b_1 _1685_ (.A(\cpu.RD_PIPELINE[3][1] ),
    .B_N(\cpu.R2_PIPELINE[1][1] ),
    .X(_0227_));
 sky130_fd_sc_hd__or2b_1 _1686_ (.A(\cpu.R2_PIPELINE[1][1] ),
    .B_N(\cpu.RD_PIPELINE[3][1] ),
    .X(_0228_));
 sky130_fd_sc_hd__o211ai_2 _1687_ (.A1(\cpu.RD_PIPELINE[3][0] ),
    .A2(_0226_),
    .B1(_0227_),
    .C1(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__xor2_1 _1688_ (.A(\cpu.RD_PIPELINE[3][2] ),
    .B(\cpu.R2_PIPELINE[1][2] ),
    .X(_0230_));
 sky130_fd_sc_hd__xor2_1 _1689_ (.A(\cpu.R2_PIPELINE[1][3] ),
    .B(\cpu.RD_PIPELINE[3][3] ),
    .X(_0231_));
 sky130_fd_sc_hd__a2111o_1 _1690_ (.A1(\cpu.RD_PIPELINE[3][0] ),
    .A2(_0226_),
    .B1(_0230_),
    .C1(_0231_),
    .D1(\cpu.RD_PIPELINE[3][4] ),
    .X(_0232_));
 sky130_fd_sc_hd__nor3_4 _1691_ (.A(_0225_),
    .B(_0229_),
    .C(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__clkbuf_4 _1692_ (.A(\cpu.INSTRUCTION_EXECUTE_3[11] ),
    .X(_0234_));
 sky130_fd_sc_hd__buf_4 _1693_ (.A(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .X(_0235_));
 sky130_fd_sc_hd__buf_4 _1694_ (.A(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .X(_0236_));
 sky130_fd_sc_hd__buf_4 _1695_ (.A(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .X(_0237_));
 sky130_fd_sc_hd__and4b_2 _1696_ (.A_N(_0234_),
    .B(_0235_),
    .C(_0236_),
    .D(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__and4b_2 _1697_ (.A_N(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .B(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .D(_0234_),
    .X(_0239_));
 sky130_fd_sc_hd__buf_4 _1698_ (.A(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _1699_ (.A1(\cpu.regFile.REGISTERS[7][1] ),
    .A2(_0238_),
    .B1(_0240_),
    .B2(\cpu.regFile.REGISTERS[11][1] ),
    .X(_0241_));
 sky130_fd_sc_hd__nor4b_4 _1700_ (.A(_0207_),
    .B(_0236_),
    .C(_0237_),
    .D_N(_0235_),
    .Y(_0242_));
 sky130_fd_sc_hd__and4bb_2 _1701_ (.A_N(_0234_),
    .B_N(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .D(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _1702_ (.A1(\cpu.regFile.REGISTERS[2][1] ),
    .A2(_0242_),
    .B1(_0243_),
    .B2(\cpu.regFile.REGISTERS[3][1] ),
    .X(_0244_));
 sky130_fd_sc_hd__or2_1 _1703_ (.A(_0241_),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__and4_2 _1704_ (.A(_0207_),
    .B(_0235_),
    .C(_0236_),
    .D(_0237_),
    .X(_0246_));
 sky130_fd_sc_hd__buf_4 _1705_ (.A(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__and4bb_2 _1706_ (.A_N(_0207_),
    .B_N(_0236_),
    .C(_0237_),
    .D(_0235_),
    .X(_0248_));
 sky130_fd_sc_hd__buf_4 _1707_ (.A(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__and4b_2 _1708_ (.A_N(_0236_),
    .B(_0237_),
    .C(_0207_),
    .D(_0235_),
    .X(_0250_));
 sky130_fd_sc_hd__and4bb_2 _1709_ (.A_N(_0236_),
    .B_N(_0237_),
    .C(_0207_),
    .D(_0235_),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _1710_ (.A1(\cpu.regFile.REGISTERS[14][1] ),
    .A2(_0250_),
    .B1(_0251_),
    .B2(\cpu.regFile.REGISTERS[10][1] ),
    .X(_0252_));
 sky130_fd_sc_hd__a221o_1 _1711_ (.A1(\cpu.regFile.REGISTERS[15][1] ),
    .A2(_0247_),
    .B1(_0249_),
    .B2(\cpu.regFile.REGISTERS[6][1] ),
    .C1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__and4bb_2 _1712_ (.A_N(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .B_N(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .D(_0234_),
    .X(_0254_));
 sky130_fd_sc_hd__nor4b_4 _1713_ (.A(_0234_),
    .B(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .D_N(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .Y(_0255_));
 sky130_fd_sc_hd__a22o_1 _1714_ (.A1(\cpu.regFile.REGISTERS[12][1] ),
    .A2(_0254_),
    .B1(_0255_),
    .B2(\cpu.regFile.REGISTERS[1][1] ),
    .X(_0256_));
 sky130_fd_sc_hd__and4bb_2 _1715_ (.A_N(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .B_N(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .D(_0234_),
    .X(_0257_));
 sky130_fd_sc_hd__and4bb_2 _1716_ (.A_N(_0234_),
    .B_N(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .D(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _1717_ (.A1(\cpu.regFile.REGISTERS[9][1] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(\cpu.regFile.REGISTERS[5][1] ),
    .X(_0259_));
 sky130_fd_sc_hd__nor4b_4 _1718_ (.A(_0234_),
    .B(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .D_N(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .Y(_0260_));
 sky130_fd_sc_hd__nor4_4 _1719_ (.A(_0207_),
    .B(_0235_),
    .C(_0236_),
    .D(_0237_),
    .Y(_0261_));
 sky130_fd_sc_hd__a21o_1 _1720_ (.A1(\cpu.regFile.REGISTERS[4][1] ),
    .A2(_0260_),
    .B1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__nor4b_4 _1721_ (.A(_0235_),
    .B(_0236_),
    .C(_0237_),
    .D_N(_0234_),
    .Y(_0263_));
 sky130_fd_sc_hd__and4b_2 _1722_ (.A_N(\cpu.INSTRUCTION_EXECUTE_3[21] ),
    .B(\cpu.INSTRUCTION_EXECUTE_3[20] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[22] ),
    .D(_0234_),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _1723_ (.A1(\cpu.regFile.REGISTERS[8][1] ),
    .A2(_0263_),
    .B1(_0264_),
    .B2(\cpu.regFile.REGISTERS[13][1] ),
    .X(_0265_));
 sky130_fd_sc_hd__or4_1 _1724_ (.A(_0256_),
    .B(_0259_),
    .C(_0262_),
    .D(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__or3_1 _1725_ (.A(_0245_),
    .B(_0253_),
    .C(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__or4_4 _1726_ (.A(_0207_),
    .B(_0235_),
    .C(_0236_),
    .D(_0237_),
    .X(_0268_));
 sky130_fd_sc_hd__or3_1 _1727_ (.A(_0225_),
    .B(_0229_),
    .C(_0232_),
    .X(_0269_));
 sky130_fd_sc_hd__buf_2 _1728_ (.A(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__o21a_1 _1729_ (.A1(\cpu.regFile.REGISTERS[0][1] ),
    .A2(_0268_),
    .B1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__inv_2 _1730_ (.A(\cpu.RD_PIPELINE[2][3] ),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _1731_ (.A(\cpu.RD_PIPELINE[2][1] ),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _1732_ (.A(\cpu.R2_PIPELINE[1][3] ),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _1733_ (.A(\cpu.R2_PIPELINE[1][1] ),
    .Y(_0275_));
 sky130_fd_sc_hd__or2_1 _1734_ (.A(\cpu.RD_PIPELINE[2][2] ),
    .B(\cpu.R2_PIPELINE[1][2] ),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_1 _1735_ (.A(\cpu.RD_PIPELINE[2][2] ),
    .B(\cpu.R2_PIPELINE[1][2] ),
    .Y(_0277_));
 sky130_fd_sc_hd__xor2_1 _1736_ (.A(\cpu.RD_PIPELINE[2][0] ),
    .B(\cpu.R2_PIPELINE[1][0] ),
    .X(_0278_));
 sky130_fd_sc_hd__a221o_1 _1737_ (.A1(\cpu.RD_PIPELINE[2][1] ),
    .A2(_0275_),
    .B1(_0276_),
    .B2(_0277_),
    .C1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__a2111o_1 _1738_ (.A1(_0274_),
    .A2(\cpu.RD_PIPELINE[2][3] ),
    .B1(\cpu.RD_PIPELINE[2][4] ),
    .C1(_0225_),
    .D1(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__a221oi_4 _1739_ (.A1(\cpu.R2_PIPELINE[1][3] ),
    .A2(_0272_),
    .B1(\cpu.R2_PIPELINE[1][1] ),
    .B2(_0273_),
    .C1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__a221oi_4 _1740_ (.A1(net160),
    .A2(_0233_),
    .B1(_0267_),
    .B2(_0271_),
    .C1(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__a221o_2 _1741_ (.A1(\cpu.R2_PIPELINE[1][3] ),
    .A2(_0272_),
    .B1(\cpu.R2_PIPELINE[1][1] ),
    .B2(_0273_),
    .C1(_0280_),
    .X(_0283_));
 sky130_fd_sc_hd__nor2_1 _1742_ (.A(net213),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__or2_1 _1743_ (.A(_0282_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__clkinv_2 _1744_ (.A(_0285_),
    .Y(\cpu.R2_DATA[1] ));
 sky130_fd_sc_hd__mux2_1 _1745_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[3] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[3] ),
    .S(_0221_),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _1746_ (.A(_0286_),
    .X(\cpu.REG_WRITE_DATA[3] ));
 sky130_fd_sc_hd__clkbuf_4 _1747_ (.A(_0281_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _1748_ (.A(net201),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__buf_4 _1749_ (.A(_0270_),
    .X(_0289_));
 sky130_fd_sc_hd__buf_6 _1750_ (.A(_0268_),
    .X(_0290_));
 sky130_fd_sc_hd__buf_4 _1751_ (.A(_0250_),
    .X(_0291_));
 sky130_fd_sc_hd__buf_4 _1752_ (.A(_0257_),
    .X(_0292_));
 sky130_fd_sc_hd__buf_4 _1753_ (.A(_0254_),
    .X(_0293_));
 sky130_fd_sc_hd__buf_4 _1754_ (.A(_0263_),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(\cpu.regFile.REGISTERS[12][3] ),
    .A2(_0293_),
    .B1(_0294_),
    .B2(\cpu.regFile.REGISTERS[8][3] ),
    .X(_0295_));
 sky130_fd_sc_hd__a221o_1 _1756_ (.A1(\cpu.regFile.REGISTERS[14][3] ),
    .A2(_0291_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][3] ),
    .C1(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__buf_4 _1757_ (.A(_0260_),
    .X(_0297_));
 sky130_fd_sc_hd__buf_4 _1758_ (.A(_0264_),
    .X(_0298_));
 sky130_fd_sc_hd__a22o_1 _1759_ (.A1(\cpu.regFile.REGISTERS[10][3] ),
    .A2(_0251_),
    .B1(_0258_),
    .B2(\cpu.regFile.REGISTERS[5][3] ),
    .X(_0299_));
 sky130_fd_sc_hd__a221o_1 _1760_ (.A1(\cpu.regFile.REGISTERS[4][3] ),
    .A2(_0297_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][3] ),
    .C1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_4 _1761_ (.A(_0238_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_4 _1762_ (.A(_0255_),
    .X(_0302_));
 sky130_fd_sc_hd__a22o_1 _1763_ (.A1(\cpu.regFile.REGISTERS[11][3] ),
    .A2(_0240_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][3] ),
    .X(_0303_));
 sky130_fd_sc_hd__a221o_1 _1764_ (.A1(\cpu.regFile.REGISTERS[7][3] ),
    .A2(_0301_),
    .B1(_0249_),
    .B2(\cpu.regFile.REGISTERS[6][3] ),
    .C1(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__buf_4 _1765_ (.A(_0242_),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _1766_ (.A1(\cpu.regFile.REGISTERS[3][3] ),
    .A2(_0243_),
    .B1(_0246_),
    .B2(\cpu.regFile.REGISTERS[15][3] ),
    .X(_0306_));
 sky130_fd_sc_hd__buf_4 _1767_ (.A(_0261_),
    .X(_0307_));
 sky130_fd_sc_hd__a211o_1 _1768_ (.A1(\cpu.regFile.REGISTERS[2][3] ),
    .A2(_0305_),
    .B1(_0306_),
    .C1(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__or3_1 _1769_ (.A(_0300_),
    .B(_0304_),
    .C(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__o22ai_4 _1770_ (.A1(\cpu.regFile.REGISTERS[0][3] ),
    .A2(_0290_),
    .B1(_0296_),
    .B2(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__nor2_1 _1771_ (.A(_0270_),
    .B(\cpu.REG_WRITE_DATA[3] ),
    .Y(_0311_));
 sky130_fd_sc_hd__a211o_2 _1772_ (.A1(_0289_),
    .A2(_0310_),
    .B1(_0311_),
    .C1(_0281_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_2 _1773_ (.A(_0288_),
    .B(_0312_),
    .Y(\cpu.R2_DATA[3] ));
 sky130_fd_sc_hd__mux2_1 _1774_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[2] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[2] ),
    .S(_0221_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _1775_ (.A(_0313_),
    .X(\cpu.REG_WRITE_DATA[2] ));
 sky130_fd_sc_hd__buf_4 _1776_ (.A(_0251_),
    .X(_0314_));
 sky130_fd_sc_hd__a22o_1 _1777_ (.A1(\cpu.regFile.REGISTERS[14][2] ),
    .A2(_0291_),
    .B1(_0314_),
    .B2(\cpu.regFile.REGISTERS[10][2] ),
    .X(_0315_));
 sky130_fd_sc_hd__a221o_1 _1778_ (.A1(\cpu.regFile.REGISTERS[15][2] ),
    .A2(_0247_),
    .B1(_0294_),
    .B2(\cpu.regFile.REGISTERS[8][2] ),
    .C1(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__buf_4 _1779_ (.A(_0258_),
    .X(_0317_));
 sky130_fd_sc_hd__a22o_1 _1780_ (.A1(\cpu.regFile.REGISTERS[9][2] ),
    .A2(_0257_),
    .B1(_0297_),
    .B2(\cpu.regFile.REGISTERS[4][2] ),
    .X(_0318_));
 sky130_fd_sc_hd__a221o_1 _1781_ (.A1(\cpu.regFile.REGISTERS[12][2] ),
    .A2(_0293_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][2] ),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_1 _1782_ (.A1(\cpu.regFile.REGISTERS[7][2] ),
    .A2(_0238_),
    .B1(_0248_),
    .B2(\cpu.regFile.REGISTERS[6][2] ),
    .X(_0320_));
 sky130_fd_sc_hd__a221o_1 _1783_ (.A1(\cpu.regFile.REGISTERS[1][2] ),
    .A2(_0302_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][2] ),
    .C1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__buf_4 _1784_ (.A(_0243_),
    .X(_0322_));
 sky130_fd_sc_hd__a22o_1 _1785_ (.A1(\cpu.regFile.REGISTERS[11][2] ),
    .A2(_0240_),
    .B1(_0322_),
    .B2(\cpu.regFile.REGISTERS[3][2] ),
    .X(_0323_));
 sky130_fd_sc_hd__a211o_1 _1786_ (.A1(\cpu.regFile.REGISTERS[2][2] ),
    .A2(_0305_),
    .B1(_0323_),
    .C1(_0307_),
    .X(_0324_));
 sky130_fd_sc_hd__or3_1 _1787_ (.A(_0319_),
    .B(_0321_),
    .C(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__o22a_2 _1788_ (.A1(\cpu.regFile.REGISTERS[0][2] ),
    .A2(_0290_),
    .B1(_0316_),
    .B2(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__o21a_1 _1789_ (.A1(_0270_),
    .A2(net155),
    .B1(_0283_),
    .X(_0327_));
 sky130_fd_sc_hd__o21ai_2 _1790_ (.A1(_0233_),
    .A2(_0326_),
    .B1(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_1 _1791_ (.A(net207),
    .B(_0287_),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_2 _1792_ (.A(_0328_),
    .B(_0329_),
    .Y(\cpu.R2_DATA[2] ));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[6] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[6] ),
    .S(_0221_),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _1794_ (.A(_0330_),
    .X(\cpu.REG_WRITE_DATA[6] ));
 sky130_fd_sc_hd__a22o_1 _1795_ (.A1(\cpu.regFile.REGISTERS[14][6] ),
    .A2(_0250_),
    .B1(_0314_),
    .B2(\cpu.regFile.REGISTERS[10][6] ),
    .X(_0331_));
 sky130_fd_sc_hd__a221o_1 _1796_ (.A1(\cpu.regFile.REGISTERS[15][6] ),
    .A2(_0247_),
    .B1(_0294_),
    .B2(\cpu.regFile.REGISTERS[8][6] ),
    .C1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_1 _1797_ (.A1(\cpu.regFile.REGISTERS[9][6] ),
    .A2(_0257_),
    .B1(_0260_),
    .B2(\cpu.regFile.REGISTERS[4][6] ),
    .X(_0333_));
 sky130_fd_sc_hd__a221o_1 _1798_ (.A1(\cpu.regFile.REGISTERS[12][6] ),
    .A2(_0254_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][6] ),
    .C1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _1799_ (.A1(\cpu.regFile.REGISTERS[1][6] ),
    .A2(_0255_),
    .B1(_0264_),
    .B2(\cpu.regFile.REGISTERS[13][6] ),
    .X(_0335_));
 sky130_fd_sc_hd__a221o_1 _1800_ (.A1(\cpu.regFile.REGISTERS[7][6] ),
    .A2(_0238_),
    .B1(_0248_),
    .B2(\cpu.regFile.REGISTERS[6][6] ),
    .C1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _1801_ (.A1(\cpu.regFile.REGISTERS[11][6] ),
    .A2(_0239_),
    .B1(_0243_),
    .B2(\cpu.regFile.REGISTERS[3][6] ),
    .X(_0337_));
 sky130_fd_sc_hd__a211o_1 _1802_ (.A1(\cpu.regFile.REGISTERS[2][6] ),
    .A2(_0242_),
    .B1(_0337_),
    .C1(_0261_),
    .X(_0338_));
 sky130_fd_sc_hd__or3_1 _1803_ (.A(_0334_),
    .B(_0336_),
    .C(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__o22a_1 _1804_ (.A1(\cpu.regFile.REGISTERS[0][6] ),
    .A2(_0268_),
    .B1(_0332_),
    .B2(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(net152),
    .A1(_0340_),
    .S(_0270_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_6 _1806_ (.A(_0283_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(net182),
    .A1(_0341_),
    .S(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_4 _1808_ (.A(_0343_),
    .X(\cpu.R2_DATA[6] ));
 sky130_fd_sc_hd__clkbuf_4 _1809_ (.A(_0221_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[5] ),
    .S(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _1811_ (.A(_0345_),
    .X(\cpu.REG_WRITE_DATA[5] ));
 sky130_fd_sc_hd__or2_1 _1812_ (.A(net189),
    .B(_0342_),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _1813_ (.A1(\cpu.regFile.REGISTERS[12][5] ),
    .A2(_0293_),
    .B1(_0263_),
    .B2(\cpu.regFile.REGISTERS[8][5] ),
    .X(_0347_));
 sky130_fd_sc_hd__a221o_1 _1814_ (.A1(\cpu.regFile.REGISTERS[14][5] ),
    .A2(_0291_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][5] ),
    .C1(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _1815_ (.A1(\cpu.regFile.REGISTERS[10][5] ),
    .A2(_0251_),
    .B1(_0258_),
    .B2(\cpu.regFile.REGISTERS[5][5] ),
    .X(_0349_));
 sky130_fd_sc_hd__a221o_1 _1816_ (.A1(\cpu.regFile.REGISTERS[4][5] ),
    .A2(_0297_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][5] ),
    .C1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _1817_ (.A1(\cpu.regFile.REGISTERS[11][5] ),
    .A2(_0239_),
    .B1(_0255_),
    .B2(\cpu.regFile.REGISTERS[1][5] ),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_1 _1818_ (.A1(\cpu.regFile.REGISTERS[7][5] ),
    .A2(_0301_),
    .B1(_0249_),
    .B2(\cpu.regFile.REGISTERS[6][5] ),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _1819_ (.A1(\cpu.regFile.REGISTERS[3][5] ),
    .A2(_0243_),
    .B1(_0246_),
    .B2(\cpu.regFile.REGISTERS[15][5] ),
    .X(_0353_));
 sky130_fd_sc_hd__a211o_1 _1820_ (.A1(\cpu.regFile.REGISTERS[2][5] ),
    .A2(_0242_),
    .B1(_0353_),
    .C1(_0261_),
    .X(_0354_));
 sky130_fd_sc_hd__or3_1 _1821_ (.A(_0350_),
    .B(_0352_),
    .C(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _1822_ (.A(_0348_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__o21a_1 _1823_ (.A1(\cpu.regFile.REGISTERS[0][5] ),
    .A2(_0268_),
    .B1(_0270_),
    .X(_0357_));
 sky130_fd_sc_hd__a221o_1 _1824_ (.A1(_0233_),
    .A2(net143),
    .B1(_0356_),
    .B2(_0357_),
    .C1(_0281_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _1825_ (.A(_0346_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_2 _1826_ (.A(_0359_),
    .X(\cpu.R2_DATA[5] ));
 sky130_fd_sc_hd__mux2_1 _1827_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[4] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[4] ),
    .S(_0221_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_2 _1828_ (.A(_0360_),
    .X(\cpu.REG_WRITE_DATA[4] ));
 sky130_fd_sc_hd__nand2_1 _1829_ (.A(net195),
    .B(_0287_),
    .Y(_0361_));
 sky130_fd_sc_hd__a22o_1 _1830_ (.A1(\cpu.regFile.REGISTERS[12][4] ),
    .A2(_0293_),
    .B1(_0294_),
    .B2(\cpu.regFile.REGISTERS[8][4] ),
    .X(_0362_));
 sky130_fd_sc_hd__a221o_1 _1831_ (.A1(\cpu.regFile.REGISTERS[14][4] ),
    .A2(_0291_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][4] ),
    .C1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _1832_ (.A1(\cpu.regFile.REGISTERS[4][4] ),
    .A2(_0297_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][4] ),
    .X(_0364_));
 sky130_fd_sc_hd__a221o_1 _1833_ (.A1(\cpu.regFile.REGISTERS[10][4] ),
    .A2(_0314_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][4] ),
    .C1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _1834_ (.A1(\cpu.regFile.REGISTERS[11][4] ),
    .A2(_0240_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][4] ),
    .X(_0366_));
 sky130_fd_sc_hd__a221o_1 _1835_ (.A1(\cpu.regFile.REGISTERS[7][4] ),
    .A2(_0301_),
    .B1(_0249_),
    .B2(\cpu.regFile.REGISTERS[6][4] ),
    .C1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__a22o_1 _1836_ (.A1(\cpu.regFile.REGISTERS[3][4] ),
    .A2(_0322_),
    .B1(_0246_),
    .B2(\cpu.regFile.REGISTERS[15][4] ),
    .X(_0368_));
 sky130_fd_sc_hd__a211o_1 _1837_ (.A1(\cpu.regFile.REGISTERS[2][4] ),
    .A2(_0305_),
    .B1(_0368_),
    .C1(_0307_),
    .X(_0369_));
 sky130_fd_sc_hd__or3_1 _1838_ (.A(_0365_),
    .B(_0367_),
    .C(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__o22ai_4 _1839_ (.A1(\cpu.regFile.REGISTERS[0][4] ),
    .A2(_0290_),
    .B1(_0363_),
    .B2(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _1840_ (.A(_0289_),
    .B(\cpu.REG_WRITE_DATA[4] ),
    .Y(_0372_));
 sky130_fd_sc_hd__a211o_2 _1841_ (.A1(_0289_),
    .A2(_0371_),
    .B1(_0372_),
    .C1(_0287_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_4 _1842_ (.A(_0361_),
    .B(_0373_),
    .Y(\cpu.R2_DATA[4] ));
 sky130_fd_sc_hd__and2_1 _1843_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[15] ),
    .B(_0344_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _1844_ (.A(_0374_),
    .X(\cpu.REG_WRITE_DATA[15] ));
 sky130_fd_sc_hd__and2_1 _1845_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[13] ),
    .B(_0344_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _1846_ (.A(_0375_),
    .X(\cpu.REG_WRITE_DATA[13] ));
 sky130_fd_sc_hd__buf_2 _1847_ (.A(_0344_),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _1848_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[12] ),
    .B(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _1849_ (.A(_0377_),
    .X(\cpu.REG_WRITE_DATA[12] ));
 sky130_fd_sc_hd__and2_1 _1850_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[11] ),
    .B(_0344_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_2 _1851_ (.A(_0378_),
    .X(\cpu.REG_WRITE_DATA[11] ));
 sky130_fd_sc_hd__and2_1 _1852_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[10] ),
    .B(_0344_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_2 _1853_ (.A(_0379_),
    .X(\cpu.REG_WRITE_DATA[10] ));
 sky130_fd_sc_hd__and2_1 _1854_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[9] ),
    .B(_0344_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _1855_ (.A(_0380_),
    .X(\cpu.REG_WRITE_DATA[9] ));
 sky130_fd_sc_hd__and2_1 _1856_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[8] ),
    .B(_0344_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _1857_ (.A(_0381_),
    .X(\cpu.REG_WRITE_DATA[8] ));
 sky130_fd_sc_hd__buf_4 _1858_ (.A(_0376_),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _1859_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[31] ),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _1860_ (.A(_0383_),
    .X(\cpu.REG_WRITE_DATA[31] ));
 sky130_fd_sc_hd__and2_1 _1861_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[30] ),
    .B(_0382_),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _1862_ (.A(_0384_),
    .X(\cpu.REG_WRITE_DATA[30] ));
 sky130_fd_sc_hd__and2_1 _1863_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[29] ),
    .B(_0382_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_2 _1864_ (.A(_0385_),
    .X(\cpu.REG_WRITE_DATA[29] ));
 sky130_fd_sc_hd__and2_1 _1865_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[28] ),
    .B(_0382_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_2 _1866_ (.A(_0386_),
    .X(\cpu.REG_WRITE_DATA[28] ));
 sky130_fd_sc_hd__and2_1 _1867_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[27] ),
    .B(_0382_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_2 _1868_ (.A(_0387_),
    .X(\cpu.REG_WRITE_DATA[27] ));
 sky130_fd_sc_hd__and2_1 _1869_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[26] ),
    .B(_0382_),
    .X(_0388_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1870_ (.A(_0388_),
    .X(\cpu.REG_WRITE_DATA[26] ));
 sky130_fd_sc_hd__and2_1 _1871_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[25] ),
    .B(_0382_),
    .X(_0389_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1872_ (.A(_0389_),
    .X(\cpu.REG_WRITE_DATA[25] ));
 sky130_fd_sc_hd__and2_1 _1873_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[24] ),
    .B(_0382_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_2 _1874_ (.A(_0390_),
    .X(\cpu.REG_WRITE_DATA[24] ));
 sky130_fd_sc_hd__and2_1 _1875_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[23] ),
    .B(_0376_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_2 _1876_ (.A(_0391_),
    .X(\cpu.REG_WRITE_DATA[23] ));
 sky130_fd_sc_hd__and2_1 _1877_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[22] ),
    .B(_0376_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_2 _1878_ (.A(_0392_),
    .X(\cpu.REG_WRITE_DATA[22] ));
 sky130_fd_sc_hd__and2_1 _1879_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[21] ),
    .B(_0344_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _1880_ (.A(_0393_),
    .X(\cpu.REG_WRITE_DATA[21] ));
 sky130_fd_sc_hd__and2_1 _1881_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[20] ),
    .B(_0376_),
    .X(_0394_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1882_ (.A(_0394_),
    .X(\cpu.REG_WRITE_DATA[20] ));
 sky130_fd_sc_hd__and2_1 _1883_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[17] ),
    .B(_0376_),
    .X(_0395_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1884_ (.A(_0395_),
    .X(\cpu.REG_WRITE_DATA[17] ));
 sky130_fd_sc_hd__and2_1 _1885_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[16] ),
    .B(_0376_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _1886_ (.A(_0396_),
    .X(\cpu.REG_WRITE_DATA[16] ));
 sky130_fd_sc_hd__xnor2_1 _1887_ (.A(\cpu.RD_PIPELINE[1][2] ),
    .B(\cpu.R2_PIPELINE[0][2] ),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _1888_ (.A(\cpu.RD_PIPELINE[1][0] ),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _1889_ (.A(\cpu.RD_PIPELINE[1][3] ),
    .Y(_0399_));
 sky130_fd_sc_hd__xnor2_1 _1890_ (.A(\cpu.RD_PIPELINE[1][1] ),
    .B(\cpu.R2_PIPELINE[0][1] ),
    .Y(_0400_));
 sky130_fd_sc_hd__o221a_1 _1891_ (.A1(_0398_),
    .A2(\cpu.R2_PIPELINE[0][0] ),
    .B1(\cpu.R2_PIPELINE[0][3] ),
    .B2(_0399_),
    .C1(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__inv_2 _1892_ (.A(\cpu.R2_PIPELINE[0][3] ),
    .Y(_0402_));
 sky130_fd_sc_hd__o31a_1 _1893_ (.A1(\cpu.R2_PIPELINE[0][1] ),
    .A2(\cpu.R2_PIPELINE[0][0] ),
    .A3(\cpu.R2_PIPELINE[0][2] ),
    .B1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_1 _1894_ (.A1(_0398_),
    .A2(\cpu.R2_PIPELINE[0][0] ),
    .B1(\cpu.R2_PIPELINE[1][3] ),
    .Y(_0404_));
 sky130_fd_sc_hd__or4_1 _1895_ (.A(\cpu.TYPE_PIPELINE[0][1] ),
    .B(\cpu.TYPE_PIPELINE[0][3] ),
    .C(\cpu.TYPE_PIPELINE[0][2] ),
    .D(\cpu.TYPE_PIPELINE[0][4] ),
    .X(_0405_));
 sky130_fd_sc_hd__o211a_1 _1896_ (.A1(\cpu.RD_PIPELINE[1][3] ),
    .A2(_0403_),
    .B1(_0404_),
    .C1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__or4b_1 _1897_ (.A(\cpu.RD_PIPELINE[1][0] ),
    .B(\cpu.RD_PIPELINE[1][3] ),
    .C(\cpu.R2_PIPELINE[1][3] ),
    .D_N(\cpu.RD_PIPELINE[1][2] ),
    .X(_0407_));
 sky130_fd_sc_hd__inv_2 _1898_ (.A(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__o2111a_1 _1899_ (.A1(\cpu.TYPE_PIPELINE[0][0] ),
    .A2(_0405_),
    .B1(_0408_),
    .C1(\cpu.RD_PIPELINE[1][1] ),
    .D1(\cpu.R1_PIPELINE[0][1] ),
    .X(_0409_));
 sky130_fd_sc_hd__a31o_1 _1900_ (.A1(_0397_),
    .A2(_0401_),
    .A3(_0406_),
    .B1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__and2_1 _1901_ (.A(\cpu.TYPE_PIPELINE[1][3] ),
    .B(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_4 _1902_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__or2b_1 _1903_ (.A(\cpu.INSTRUCTION_DECODE_2[11] ),
    .B_N(\cpu.INSTRUCTION_DECODE_2[0] ),
    .X(_0413_));
 sky130_fd_sc_hd__a21oi_1 _1904_ (.A1(\cpu.TYPE_PIPELINE[1][4] ),
    .A2(_0413_),
    .B1(_0213_),
    .Y(_0414_));
 sky130_fd_sc_hd__nor2_1 _1905_ (.A(_0412_),
    .B(_0414_),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_1 _1906_ (.A(\cpu.TYPE_PIPELINE[1][3] ),
    .B(_0410_),
    .Y(_0415_));
 sky130_fd_sc_hd__buf_4 _1907_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__and3b_1 _1908_ (.A_N(_0213_),
    .B(_0416_),
    .C(_0413_),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _1909_ (.A(\cpu.INSTRUCTION_DECODE_2[5] ),
    .B(_0415_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1910_ (.A(_0418_),
    .X(_0120_));
 sky130_fd_sc_hd__and2b_1 _1911_ (.A_N(_0413_),
    .B(_0120_),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _1912_ (.A1(\cpu.TYPE_PIPELINE[1][2] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(_0212_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_2 _1913_ (.A(_0416_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _1914_ (.A(\cpu.INSTRUCTION_DECODE_2[5] ),
    .B(_0413_),
    .Y(_0421_));
 sky130_fd_sc_hd__a32o_1 _1915_ (.A1(_0212_),
    .A2(_0420_),
    .A3(_0421_),
    .B1(_0417_),
    .B2(\cpu.TYPE_PIPELINE[1][3] ),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_1 _1916_ (.A1(\cpu.TYPE_PIPELINE[1][1] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(\cpu.INSTRUCTION_DECODE_2[4] ),
    .X(_0006_));
 sky130_fd_sc_hd__nand3b_4 _1917_ (.A_N(\cpu.INSTRUCTION_WRITEBACK_5[11] ),
    .B(\cpu.INSTRUCTION_WRITEBACK_5[4] ),
    .C(\cpu.INSTRUCTION_WRITEBACK_5[0] ),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _1918_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[8] ),
    .Y(_0423_));
 sky130_fd_sc_hd__a211o_1 _1919_ (.A1(_0382_),
    .A2(_0422_),
    .B1(\cpu.INSTRUCTION_WRITEBACK_5[7] ),
    .C1(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_2 _1920_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[9] ),
    .X(_0425_));
 sky130_fd_sc_hd__buf_2 _1921_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[10] ),
    .X(_0426_));
 sky130_fd_sc_hd__or3b_1 _1922_ (.A(_0424_),
    .B(_0425_),
    .C_N(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__buf_2 _1923_ (.A(_0427_),
    .X(_0023_));
 sky130_fd_sc_hd__clkinv_2 _1924_ (.A(_0344_),
    .Y(_0428_));
 sky130_fd_sc_hd__and3b_1 _1925_ (.A_N(\cpu.INSTRUCTION_WRITEBACK_5[11] ),
    .B(\cpu.INSTRUCTION_WRITEBACK_5[4] ),
    .C(\cpu.INSTRUCTION_WRITEBACK_5[0] ),
    .X(_0429_));
 sky130_fd_sc_hd__o211a_1 _1926_ (.A1(_0428_),
    .A2(_0429_),
    .B1(\cpu.INSTRUCTION_WRITEBACK_5[7] ),
    .C1(\cpu.INSTRUCTION_WRITEBACK_5[8] ),
    .X(_0430_));
 sky130_fd_sc_hd__nand3_1 _1927_ (.A(_0425_),
    .B(_0426_),
    .C(_0430_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand3b_4 _1928_ (.A_N(_0425_),
    .B(_0426_),
    .C(_0430_),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2_1 _1929_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[9] ),
    .B(\cpu.INSTRUCTION_WRITEBACK_5[10] ),
    .Y(_0431_));
 sky130_fd_sc_hd__a211o_1 _1930_ (.A1(_0382_),
    .A2(_0422_),
    .B1(\cpu.INSTRUCTION_WRITEBACK_5[7] ),
    .C1(\cpu.INSTRUCTION_WRITEBACK_5[8] ),
    .X(_0432_));
 sky130_fd_sc_hd__or2_1 _1931_ (.A(_0431_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_2 _1932_ (.A(_0433_),
    .X(_0025_));
 sky130_fd_sc_hd__o211ai_2 _1933_ (.A1(_0428_),
    .A2(_0429_),
    .B1(\cpu.INSTRUCTION_WRITEBACK_5[7] ),
    .C1(_0423_),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_1 _1934_ (.A(_0431_),
    .B(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _1935_ (.A(_0435_),
    .X(_0026_));
 sky130_fd_sc_hd__or3_1 _1936_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[9] ),
    .B(\cpu.INSTRUCTION_WRITEBACK_5[10] ),
    .C(_0434_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1937_ (.A(_0436_),
    .X(_0014_));
 sky130_fd_sc_hd__or3_1 _1938_ (.A(\cpu.INSTRUCTION_WRITEBACK_5[9] ),
    .B(\cpu.INSTRUCTION_WRITEBACK_5[10] ),
    .C(_0424_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1939_ (.A(_0437_),
    .X(_0015_));
 sky130_fd_sc_hd__or3b_1 _1940_ (.A(_0425_),
    .B(_0426_),
    .C_N(_0430_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _1941_ (.A(_0438_),
    .X(_0016_));
 sky130_fd_sc_hd__or3b_1 _1942_ (.A(_0426_),
    .B(_0432_),
    .C_N(_0425_),
    .X(_0439_));
 sky130_fd_sc_hd__buf_2 _1943_ (.A(_0439_),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _1944_ (.A(_0424_),
    .B(_0431_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_4 _1945_ (.A(_0440_),
    .X(_0027_));
 sky130_fd_sc_hd__or3b_1 _1946_ (.A(_0426_),
    .B(_0434_),
    .C_N(_0425_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _1947_ (.A(_0441_),
    .X(_0018_));
 sky130_fd_sc_hd__or3b_1 _1948_ (.A(_0426_),
    .B(_0424_),
    .C_N(_0425_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _1949_ (.A(_0442_),
    .X(_0019_));
 sky130_fd_sc_hd__nand3b_1 _1950_ (.A_N(_0426_),
    .B(_0430_),
    .C(_0425_),
    .Y(_0020_));
 sky130_fd_sc_hd__or3b_1 _1951_ (.A(_0432_),
    .B(_0425_),
    .C_N(_0426_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _1952_ (.A(_0443_),
    .X(_0021_));
 sky130_fd_sc_hd__or3b_1 _1953_ (.A(_0434_),
    .B(_0425_),
    .C_N(_0426_),
    .X(_0444_));
 sky130_fd_sc_hd__buf_2 _1954_ (.A(_0444_),
    .X(_0022_));
 sky130_fd_sc_hd__a221o_1 _1955_ (.A1(\cpu.TYPE_PIPELINE[1][0] ),
    .A2(_0417_),
    .B1(_0421_),
    .B2(\cpu.INSTRUCTION_DECODE_2[4] ),
    .C1(_0412_),
    .X(_0005_));
 sky130_fd_sc_hd__or2b_1 _1956_ (.A(\cpu.PC[2] ),
    .B_N(\cpu.PC[5] ),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_2 _1957_ (.A(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _1958_ (.A1(_0218_),
    .A2(_0446_),
    .B1(_0215_),
    .X(_0000_));
 sky130_fd_sc_hd__nor2_2 _1959_ (.A(_0215_),
    .B(_0446_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_1 _1960_ (.A(_0219_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _1961_ (.A(_0000_),
    .B(_0447_),
    .Y(_0003_));
 sky130_fd_sc_hd__or4bb_2 _1962_ (.A(\cpu.INSTRUCTION_MEMORY_4[4] ),
    .B(\cpu.INSTRUCTION_MEMORY_4[11] ),
    .C_N(\cpu.INSTRUCTION_MEMORY_4[0] ),
    .D_N(\cpu.INSTRUCTION_MEMORY_4[5] ),
    .X(_0448_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1963_ (.A(_0448_),
    .X(_0010_));
 sky130_fd_sc_hd__inv_2 _1964_ (.A(\cpu.immediateExtractor.VALUE[31] ),
    .Y(_0449_));
 sky130_fd_sc_hd__buf_6 _1965_ (.A(_0342_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_8 _1966_ (.A(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_1 _1967_ (.A(_0428_),
    .B(_0289_),
    .Y(_0452_));
 sky130_fd_sc_hd__buf_2 _1968_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__buf_2 _1969_ (.A(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_4 _1970_ (.A(_0290_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_4 _1971_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__buf_4 _1972_ (.A(_0305_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _1973_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_4 _1974_ (.A(_0314_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_4 _1975_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__buf_4 _1976_ (.A(_0240_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_4 _1977_ (.A(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_4 _1978_ (.A(_0249_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_4 _1979_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _1980_ (.A1(\cpu.regFile.REGISTERS[11][31] ),
    .A2(_0462_),
    .B1(_0464_),
    .B2(\cpu.regFile.REGISTERS[6][31] ),
    .X(_0465_));
 sky130_fd_sc_hd__a221o_1 _1981_ (.A1(\cpu.regFile.REGISTERS[2][31] ),
    .A2(_0458_),
    .B1(_0460_),
    .B2(\cpu.regFile.REGISTERS[10][31] ),
    .C1(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__buf_4 _1982_ (.A(_0301_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_4 _1983_ (.A(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_4 _1984_ (.A(_0247_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_4 _1985_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_4 _1986_ (.A(_0322_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_4 _1987_ (.A(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__buf_4 _1988_ (.A(_0291_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_4 _1989_ (.A(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _1990_ (.A1(\cpu.regFile.REGISTERS[3][31] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][31] ),
    .X(_0475_));
 sky130_fd_sc_hd__a221o_1 _1991_ (.A1(\cpu.regFile.REGISTERS[7][31] ),
    .A2(_0468_),
    .B1(_0470_),
    .B2(\cpu.regFile.REGISTERS[15][31] ),
    .C1(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__buf_4 _1992_ (.A(_0292_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_4 _1993_ (.A(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_4 _1994_ (.A(_0294_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_4 _1995_ (.A(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_4 _1996_ (.A(_0317_),
    .X(_0481_));
 sky130_fd_sc_hd__buf_4 _1997_ (.A(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_4 _1998_ (.A(_0298_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_4 _1999_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a22o_1 _2000_ (.A1(\cpu.regFile.REGISTERS[5][31] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][31] ),
    .X(_0485_));
 sky130_fd_sc_hd__a221o_1 _2001_ (.A1(\cpu.regFile.REGISTERS[9][31] ),
    .A2(_0478_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][31] ),
    .C1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_4 _2002_ (.A(_0302_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_4 _2003_ (.A(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__buf_4 _2004_ (.A(_0293_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_4 _2005_ (.A(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_4 _2006_ (.A(_0297_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_4 _2007_ (.A(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__a22o_1 _2008_ (.A1(\cpu.regFile.REGISTERS[12][31] ),
    .A2(_0490_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][31] ),
    .X(_0493_));
 sky130_fd_sc_hd__buf_4 _2009_ (.A(_0307_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_4 _2010_ (.A(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__a211o_1 _2011_ (.A1(\cpu.regFile.REGISTERS[1][31] ),
    .A2(_0488_),
    .B1(_0493_),
    .C1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__or3_1 _2012_ (.A(_0476_),
    .B(_0486_),
    .C(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_4 _2013_ (.A(_0289_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _2014_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__o221a_1 _2015_ (.A1(\cpu.regFile.REGISTERS[0][31] ),
    .A2(_0456_),
    .B1(_0466_),
    .B2(_0497_),
    .C1(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__buf_2 _2016_ (.A(_0287_),
    .X(_0501_));
 sky130_fd_sc_hd__buf_2 _2017_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a211o_1 _2018_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[31] ),
    .A2(_0454_),
    .B1(_0500_),
    .C1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o21ai_4 _2019_ (.A1(\cpu.ALU_OUT_MEMORY_4[31] ),
    .A2(_0451_),
    .B1(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__a21oi_1 _2020_ (.A1(\cpu.INSTRUCTION_EXECUTE_3[4] ),
    .A2(\cpu.INSTRUCTION_EXECUTE_3[5] ),
    .B1(_0207_),
    .Y(_0505_));
 sky130_fd_sc_hd__a21o_2 _2021_ (.A1(\cpu.INSTRUCTION_EXECUTE_3[0] ),
    .A2(_0505_),
    .B1(_0209_),
    .X(_0506_));
 sky130_fd_sc_hd__inv_2 _2022_ (.A(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__clkbuf_2 _2023_ (.A(_0507_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2024_ (.A0(_0449_),
    .A1(_0504_),
    .S(net126),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_4 _2025_ (.A(_0211_),
    .X(_0509_));
 sky130_fd_sc_hd__buf_4 _2026_ (.A(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_4 _2027_ (.A(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__buf_4 _2028_ (.A(\cpu.INSTRUCTION_EXECUTE_3[16] ),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_4 _2029_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_4 _2030_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _2031_ (.A0(\cpu.regFile.REGISTERS[0][31] ),
    .A1(\cpu.regFile.REGISTERS[6][31] ),
    .S(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__inv_2 _2032_ (.A(\cpu.R1_PIPELINE[1][1] ),
    .Y(_0516_));
 sky130_fd_sc_hd__nor2_1 _2033_ (.A(\cpu.TYPE_PIPELINE[1][0] ),
    .B(_0223_),
    .Y(_0517_));
 sky130_fd_sc_hd__or4b_1 _2034_ (.A(\cpu.RD_PIPELINE[3][0] ),
    .B(\cpu.RD_PIPELINE[3][3] ),
    .C(\cpu.RD_PIPELINE[3][4] ),
    .D_N(\cpu.RD_PIPELINE[3][2] ),
    .X(_0518_));
 sky130_fd_sc_hd__or4b_4 _2035_ (.A(_0516_),
    .B(_0517_),
    .C(_0518_),
    .D_N(\cpu.RD_PIPELINE[3][1] ),
    .X(_0519_));
 sky130_fd_sc_hd__buf_4 _2036_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_4 _2037_ (.A(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_4 _2038_ (.A(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(net95),
    .A1(_0515_),
    .S(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__or4b_1 _2040_ (.A(\cpu.RD_PIPELINE[2][0] ),
    .B(\cpu.RD_PIPELINE[2][3] ),
    .C(\cpu.RD_PIPELINE[2][4] ),
    .D_N(\cpu.RD_PIPELINE[2][2] ),
    .X(_0524_));
 sky130_fd_sc_hd__or4_4 _2041_ (.A(_0516_),
    .B(_0273_),
    .C(_0517_),
    .D(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_4 _2042_ (.A(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_4 _2043_ (.A(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_4 _2044_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_2 _2045_ (.A0(\cpu.ALU_OUT_MEMORY_4[31] ),
    .A1(_0523_),
    .S(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__nand2_1 _2046_ (.A(_0511_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__or2b_1 _2047_ (.A(_0508_),
    .B_N(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _2048_ (.A0(\cpu.regFile.REGISTERS[0][25] ),
    .A1(\cpu.regFile.REGISTERS[6][25] ),
    .S(_0514_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _2049_ (.A0(net82),
    .A1(_0532_),
    .S(_0522_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_2 _2050_ (.A0(\cpu.ALU_OUT_MEMORY_4[25] ),
    .A1(_0533_),
    .S(_0528_),
    .X(_0534_));
 sky130_fd_sc_hd__and2_1 _2051_ (.A(_0511_),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_4 _2052_ (.A(_0506_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_4 _2053_ (.A(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _2054_ (.A1(\cpu.regFile.REGISTERS[5][25] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][25] ),
    .X(_0538_));
 sky130_fd_sc_hd__a221o_1 _2055_ (.A1(\cpu.regFile.REGISTERS[11][25] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][25] ),
    .C1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__a22o_1 _2056_ (.A1(\cpu.regFile.REGISTERS[7][25] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][25] ),
    .X(_0540_));
 sky130_fd_sc_hd__a221o_1 _2057_ (.A1(\cpu.regFile.REGISTERS[15][25] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][25] ),
    .C1(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__a22o_1 _2058_ (.A1(\cpu.regFile.REGISTERS[2][25] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][25] ),
    .X(_0542_));
 sky130_fd_sc_hd__a221o_1 _2059_ (.A1(\cpu.regFile.REGISTERS[3][25] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][25] ),
    .C1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _2060_ (.A1(\cpu.regFile.REGISTERS[10][25] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][25] ),
    .X(_0544_));
 sky130_fd_sc_hd__a211o_1 _2061_ (.A1(\cpu.regFile.REGISTERS[6][25] ),
    .A2(_0464_),
    .B1(_0544_),
    .C1(_0495_),
    .X(_0545_));
 sky130_fd_sc_hd__or3_1 _2062_ (.A(_0541_),
    .B(_0543_),
    .C(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__o221a_1 _2063_ (.A1(\cpu.regFile.REGISTERS[0][25] ),
    .A2(_0456_),
    .B1(_0539_),
    .B2(_0546_),
    .C1(_0499_),
    .X(_0547_));
 sky130_fd_sc_hd__a211o_1 _2064_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[25] ),
    .A2(_0454_),
    .B1(_0547_),
    .C1(_0502_),
    .X(_0548_));
 sky130_fd_sc_hd__o21ai_4 _2065_ (.A1(\cpu.ALU_OUT_MEMORY_4[25] ),
    .A2(_0451_),
    .B1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_2 _2066_ (.A(\cpu.immediateExtractor.VALUE[10] ),
    .B(_0506_),
    .Y(_0550_));
 sky130_fd_sc_hd__buf_4 _2067_ (.A(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__o21ai_1 _2068_ (.A1(_0537_),
    .A2(_0549_),
    .B1(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _2069_ (.A(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__mux2_1 _2070_ (.A0(\cpu.regFile.REGISTERS[0][26] ),
    .A1(\cpu.regFile.REGISTERS[6][26] ),
    .S(_0514_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _2071_ (.A0(net84),
    .A1(_0554_),
    .S(_0522_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(\cpu.ALU_OUT_MEMORY_4[26] ),
    .A1(_0555_),
    .S(_0528_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _2073_ (.A(_0510_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a22o_1 _2074_ (.A1(\cpu.regFile.REGISTERS[5][26] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][26] ),
    .X(_0558_));
 sky130_fd_sc_hd__a221o_1 _2075_ (.A1(\cpu.regFile.REGISTERS[11][26] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][26] ),
    .C1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _2076_ (.A1(\cpu.regFile.REGISTERS[7][26] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][26] ),
    .X(_0560_));
 sky130_fd_sc_hd__a221o_1 _2077_ (.A1(\cpu.regFile.REGISTERS[15][26] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][26] ),
    .C1(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_1 _2078_ (.A1(\cpu.regFile.REGISTERS[2][26] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][26] ),
    .X(_0562_));
 sky130_fd_sc_hd__a221o_1 _2079_ (.A1(\cpu.regFile.REGISTERS[3][26] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][26] ),
    .C1(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _2080_ (.A1(\cpu.regFile.REGISTERS[10][26] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][26] ),
    .X(_0564_));
 sky130_fd_sc_hd__a211o_1 _2081_ (.A1(\cpu.regFile.REGISTERS[6][26] ),
    .A2(_0464_),
    .B1(_0564_),
    .C1(_0495_),
    .X(_0565_));
 sky130_fd_sc_hd__or3_1 _2082_ (.A(_0561_),
    .B(_0563_),
    .C(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__o221a_1 _2083_ (.A1(\cpu.regFile.REGISTERS[0][26] ),
    .A2(_0456_),
    .B1(_0559_),
    .B2(_0566_),
    .C1(_0499_),
    .X(_0567_));
 sky130_fd_sc_hd__a211o_1 _2084_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[26] ),
    .A2(_0454_),
    .B1(_0567_),
    .C1(_0502_),
    .X(_0568_));
 sky130_fd_sc_hd__o21ai_4 _2085_ (.A1(\cpu.ALU_OUT_MEMORY_4[26] ),
    .A2(_0451_),
    .B1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__o21ai_2 _2086_ (.A1(_0537_),
    .A2(_0569_),
    .B1(_0551_),
    .Y(_0570_));
 sky130_fd_sc_hd__mux2_1 _2087_ (.A0(\cpu.regFile.REGISTERS[0][27] ),
    .A1(\cpu.regFile.REGISTERS[6][27] ),
    .S(_0514_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _2088_ (.A0(net86),
    .A1(_0571_),
    .S(_0522_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _2089_ (.A0(\cpu.ALU_OUT_MEMORY_4[27] ),
    .A1(_0572_),
    .S(_0528_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _2090_ (.A(_0510_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__and2_1 _2091_ (.A(\cpu.immediateExtractor.VALUE[10] ),
    .B(_0506_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_4 _2092_ (.A(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _2093_ (.A1(\cpu.regFile.REGISTERS[5][27] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][27] ),
    .X(_0577_));
 sky130_fd_sc_hd__a221o_1 _2094_ (.A1(\cpu.regFile.REGISTERS[11][27] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][27] ),
    .C1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__a22o_1 _2095_ (.A1(\cpu.regFile.REGISTERS[7][27] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][27] ),
    .X(_0579_));
 sky130_fd_sc_hd__a221o_1 _2096_ (.A1(\cpu.regFile.REGISTERS[15][27] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][27] ),
    .C1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _2097_ (.A1(\cpu.regFile.REGISTERS[2][27] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][27] ),
    .X(_0581_));
 sky130_fd_sc_hd__a221o_1 _2098_ (.A1(\cpu.regFile.REGISTERS[3][27] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][27] ),
    .C1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__a22o_1 _2099_ (.A1(\cpu.regFile.REGISTERS[10][27] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][27] ),
    .X(_0583_));
 sky130_fd_sc_hd__a211o_1 _2100_ (.A1(\cpu.regFile.REGISTERS[6][27] ),
    .A2(_0464_),
    .B1(_0583_),
    .C1(_0495_),
    .X(_0584_));
 sky130_fd_sc_hd__or3_2 _2101_ (.A(_0580_),
    .B(_0582_),
    .C(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__o221a_1 _2102_ (.A1(\cpu.regFile.REGISTERS[0][27] ),
    .A2(_0456_),
    .B1(_0578_),
    .B2(_0585_),
    .C1(_0499_),
    .X(_0586_));
 sky130_fd_sc_hd__a211o_1 _2103_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[27] ),
    .A2(_0454_),
    .B1(_0586_),
    .C1(_0502_),
    .X(_0587_));
 sky130_fd_sc_hd__o21ai_4 _2104_ (.A1(\cpu.ALU_OUT_MEMORY_4[27] ),
    .A2(_0451_),
    .B1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__nor2_1 _2105_ (.A(_0537_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _2106_ (.A(_0576_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _2107_ (.A(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__a22oi_1 _2108_ (.A1(_0557_),
    .A2(_0570_),
    .B1(_0574_),
    .B2(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__o21ai_1 _2109_ (.A1(_0557_),
    .A2(_0570_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__nor2_1 _2110_ (.A(_0574_),
    .B(_0591_),
    .Y(_0594_));
 sky130_fd_sc_hd__a211o_1 _2111_ (.A1(_0535_),
    .A2(_0553_),
    .B1(_0593_),
    .C1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _2112_ (.A0(\cpu.regFile.REGISTERS[0][29] ),
    .A1(\cpu.regFile.REGISTERS[6][29] ),
    .S(_0514_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _2113_ (.A0(net90),
    .A1(_0596_),
    .S(_0522_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_2 _2114_ (.A0(\cpu.ALU_OUT_MEMORY_4[29] ),
    .A1(_0597_),
    .S(_0528_),
    .X(_0598_));
 sky130_fd_sc_hd__nand2_1 _2115_ (.A(_0511_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__inv_2 _2116_ (.A(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__a22o_1 _2117_ (.A1(\cpu.regFile.REGISTERS[5][29] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][29] ),
    .X(_0601_));
 sky130_fd_sc_hd__a221o_1 _2118_ (.A1(\cpu.regFile.REGISTERS[11][29] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][29] ),
    .C1(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _2119_ (.A1(\cpu.regFile.REGISTERS[7][29] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][29] ),
    .X(_0603_));
 sky130_fd_sc_hd__a221o_1 _2120_ (.A1(\cpu.regFile.REGISTERS[15][29] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][29] ),
    .C1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__a22o_1 _2121_ (.A1(\cpu.regFile.REGISTERS[2][29] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][29] ),
    .X(_0605_));
 sky130_fd_sc_hd__a221o_1 _2122_ (.A1(\cpu.regFile.REGISTERS[3][29] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][29] ),
    .C1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__a22o_1 _2123_ (.A1(\cpu.regFile.REGISTERS[10][29] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][29] ),
    .X(_0607_));
 sky130_fd_sc_hd__a211o_1 _2124_ (.A1(\cpu.regFile.REGISTERS[6][29] ),
    .A2(_0464_),
    .B1(_0607_),
    .C1(_0495_),
    .X(_0608_));
 sky130_fd_sc_hd__or3_1 _2125_ (.A(_0604_),
    .B(_0606_),
    .C(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__o221a_1 _2126_ (.A1(\cpu.regFile.REGISTERS[0][29] ),
    .A2(_0456_),
    .B1(_0602_),
    .B2(_0609_),
    .C1(_0499_),
    .X(_0610_));
 sky130_fd_sc_hd__a211o_1 _2127_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[29] ),
    .A2(_0454_),
    .B1(_0610_),
    .C1(_0502_),
    .X(_0611_));
 sky130_fd_sc_hd__o21ai_4 _2128_ (.A1(\cpu.ALU_OUT_MEMORY_4[29] ),
    .A2(_0451_),
    .B1(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__or2_1 _2129_ (.A(_0537_),
    .B(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__and2_1 _2130_ (.A(_0551_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _2131_ (.A0(\cpu.regFile.REGISTERS[0][28] ),
    .A1(\cpu.regFile.REGISTERS[6][28] ),
    .S(_0514_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _2132_ (.A0(net88),
    .A1(_0615_),
    .S(_0522_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _2133_ (.A0(\cpu.ALU_OUT_MEMORY_4[28] ),
    .A1(_0616_),
    .S(_0528_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2_1 _2134_ (.A(_0511_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__a22o_1 _2135_ (.A1(\cpu.regFile.REGISTERS[5][28] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][28] ),
    .X(_0619_));
 sky130_fd_sc_hd__a221o_1 _2136_ (.A1(\cpu.regFile.REGISTERS[11][28] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][28] ),
    .C1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _2137_ (.A1(\cpu.regFile.REGISTERS[7][28] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][28] ),
    .X(_0621_));
 sky130_fd_sc_hd__a221o_1 _2138_ (.A1(\cpu.regFile.REGISTERS[15][28] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][28] ),
    .C1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _2139_ (.A1(\cpu.regFile.REGISTERS[3][28] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][28] ),
    .X(_0623_));
 sky130_fd_sc_hd__a221o_1 _2140_ (.A1(\cpu.regFile.REGISTERS[2][28] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][28] ),
    .C1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__a22o_1 _2141_ (.A1(\cpu.regFile.REGISTERS[10][28] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][28] ),
    .X(_0625_));
 sky130_fd_sc_hd__a211o_1 _2142_ (.A1(\cpu.regFile.REGISTERS[6][28] ),
    .A2(_0464_),
    .B1(_0625_),
    .C1(_0495_),
    .X(_0626_));
 sky130_fd_sc_hd__or3_1 _2143_ (.A(_0622_),
    .B(_0624_),
    .C(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__o221a_1 _2144_ (.A1(\cpu.regFile.REGISTERS[0][28] ),
    .A2(_0456_),
    .B1(_0620_),
    .B2(_0627_),
    .C1(_0499_),
    .X(_0628_));
 sky130_fd_sc_hd__a211o_1 _2145_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[28] ),
    .A2(_0454_),
    .B1(_0628_),
    .C1(_0502_),
    .X(_0629_));
 sky130_fd_sc_hd__o21ai_4 _2146_ (.A1(\cpu.ALU_OUT_MEMORY_4[28] ),
    .A2(_0451_),
    .B1(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__o21ai_2 _2147_ (.A1(_0537_),
    .A2(_0630_),
    .B1(_0551_),
    .Y(_0631_));
 sky130_fd_sc_hd__a2bb2o_1 _2148_ (.A1_N(_0600_),
    .A2_N(_0614_),
    .B1(_0618_),
    .B2(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__nor2_1 _2149_ (.A(_0618_),
    .B(_0631_),
    .Y(_0633_));
 sky130_fd_sc_hd__mux2_1 _2150_ (.A0(\cpu.regFile.REGISTERS[0][24] ),
    .A1(\cpu.regFile.REGISTERS[6][24] ),
    .S(_0514_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _2151_ (.A0(net80),
    .A1(_0634_),
    .S(_0522_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _2152_ (.A0(\cpu.ALU_OUT_MEMORY_4[24] ),
    .A1(_0635_),
    .S(_0528_),
    .X(_0636_));
 sky130_fd_sc_hd__and2_1 _2153_ (.A(_0510_),
    .B(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__a22o_1 _2154_ (.A1(\cpu.regFile.REGISTERS[5][24] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][24] ),
    .X(_0638_));
 sky130_fd_sc_hd__a221o_1 _2155_ (.A1(\cpu.regFile.REGISTERS[11][24] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][24] ),
    .C1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _2156_ (.A1(\cpu.regFile.REGISTERS[7][24] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][24] ),
    .X(_0640_));
 sky130_fd_sc_hd__a221o_1 _2157_ (.A1(\cpu.regFile.REGISTERS[15][24] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][24] ),
    .C1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__a22o_1 _2158_ (.A1(\cpu.regFile.REGISTERS[2][24] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][24] ),
    .X(_0642_));
 sky130_fd_sc_hd__a221o_1 _2159_ (.A1(\cpu.regFile.REGISTERS[3][24] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][24] ),
    .C1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a22o_1 _2160_ (.A1(\cpu.regFile.REGISTERS[10][24] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][24] ),
    .X(_0644_));
 sky130_fd_sc_hd__a211o_1 _2161_ (.A1(\cpu.regFile.REGISTERS[6][24] ),
    .A2(_0464_),
    .B1(_0644_),
    .C1(_0495_),
    .X(_0645_));
 sky130_fd_sc_hd__or3_1 _2162_ (.A(_0641_),
    .B(_0643_),
    .C(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__o221a_1 _2163_ (.A1(\cpu.regFile.REGISTERS[0][24] ),
    .A2(_0456_),
    .B1(_0639_),
    .B2(_0646_),
    .C1(_0499_),
    .X(_0647_));
 sky130_fd_sc_hd__a211o_1 _2164_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[24] ),
    .A2(_0454_),
    .B1(_0647_),
    .C1(_0502_),
    .X(_0648_));
 sky130_fd_sc_hd__o21ai_4 _2165_ (.A1(\cpu.ALU_OUT_MEMORY_4[24] ),
    .A2(_0451_),
    .B1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nor2_1 _2166_ (.A(_0537_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _2167_ (.A(_0576_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__and2_1 _2168_ (.A(_0637_),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__o22a_1 _2169_ (.A1(_0535_),
    .A2(_0553_),
    .B1(_0637_),
    .B2(_0651_),
    .X(_0653_));
 sky130_fd_sc_hd__or3b_1 _2170_ (.A(_0633_),
    .B(_0652_),
    .C_N(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _2171_ (.A0(\cpu.regFile.REGISTERS[0][30] ),
    .A1(\cpu.regFile.REGISTERS[6][30] ),
    .S(_0514_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _2172_ (.A0(net93),
    .A1(_0655_),
    .S(_0522_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_2 _2173_ (.A0(\cpu.ALU_OUT_MEMORY_4[30] ),
    .A1(_0656_),
    .S(_0528_),
    .X(_0657_));
 sky130_fd_sc_hd__and2_1 _2174_ (.A(_0511_),
    .B(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__a22o_1 _2175_ (.A1(\cpu.regFile.REGISTERS[5][30] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][30] ),
    .X(_0659_));
 sky130_fd_sc_hd__a221o_1 _2176_ (.A1(\cpu.regFile.REGISTERS[11][30] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][30] ),
    .C1(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _2177_ (.A1(\cpu.regFile.REGISTERS[7][30] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][30] ),
    .X(_0661_));
 sky130_fd_sc_hd__a221o_1 _2178_ (.A1(\cpu.regFile.REGISTERS[15][30] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][30] ),
    .C1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__a22o_1 _2179_ (.A1(\cpu.regFile.REGISTERS[2][30] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][30] ),
    .X(_0663_));
 sky130_fd_sc_hd__a221o_1 _2180_ (.A1(\cpu.regFile.REGISTERS[3][30] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][30] ),
    .C1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__a22o_1 _2181_ (.A1(\cpu.regFile.REGISTERS[10][30] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][30] ),
    .X(_0665_));
 sky130_fd_sc_hd__a211o_1 _2182_ (.A1(\cpu.regFile.REGISTERS[6][30] ),
    .A2(_0464_),
    .B1(_0665_),
    .C1(_0495_),
    .X(_0666_));
 sky130_fd_sc_hd__or3_1 _2183_ (.A(_0662_),
    .B(_0664_),
    .C(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__o221a_1 _2184_ (.A1(\cpu.regFile.REGISTERS[0][30] ),
    .A2(_0456_),
    .B1(_0660_),
    .B2(_0667_),
    .C1(_0499_),
    .X(_0668_));
 sky130_fd_sc_hd__a211o_1 _2185_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[30] ),
    .A2(_0454_),
    .B1(_0668_),
    .C1(_0502_),
    .X(_0669_));
 sky130_fd_sc_hd__o21ai_4 _2186_ (.A1(\cpu.ALU_OUT_MEMORY_4[30] ),
    .A2(_0451_),
    .B1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__o21a_1 _2187_ (.A1(_0537_),
    .A2(_0670_),
    .B1(_0551_),
    .X(_0671_));
 sky130_fd_sc_hd__xnor2_1 _2188_ (.A(_0530_),
    .B(_0508_),
    .Y(_0672_));
 sky130_fd_sc_hd__o21ai_1 _2189_ (.A1(_0658_),
    .A2(_0671_),
    .B1(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__a221o_1 _2190_ (.A1(_0658_),
    .A2(_0671_),
    .B1(_0600_),
    .B2(_0614_),
    .C1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__or4_1 _2191_ (.A(_0595_),
    .B(_0632_),
    .C(_0654_),
    .D(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _2192_ (.A0(\cpu.regFile.REGISTERS[0][22] ),
    .A1(\cpu.regFile.REGISTERS[6][22] ),
    .S(_0514_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _2193_ (.A0(net119),
    .A1(_0676_),
    .S(_0522_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_2 _2194_ (.A0(\cpu.ALU_OUT_MEMORY_4[22] ),
    .A1(_0677_),
    .S(_0528_),
    .X(_0678_));
 sky130_fd_sc_hd__nand2_2 _2195_ (.A(_0510_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__a22o_1 _2196_ (.A1(\cpu.regFile.REGISTERS[5][22] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][22] ),
    .X(_0680_));
 sky130_fd_sc_hd__a221o_1 _2197_ (.A1(\cpu.regFile.REGISTERS[11][22] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][22] ),
    .C1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__a22o_1 _2198_ (.A1(\cpu.regFile.REGISTERS[7][22] ),
    .A2(_0467_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][22] ),
    .X(_0682_));
 sky130_fd_sc_hd__a221o_1 _2199_ (.A1(\cpu.regFile.REGISTERS[15][22] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][22] ),
    .C1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__a22o_1 _2200_ (.A1(\cpu.regFile.REGISTERS[2][22] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][22] ),
    .X(_0684_));
 sky130_fd_sc_hd__a221o_1 _2201_ (.A1(\cpu.regFile.REGISTERS[3][22] ),
    .A2(_0471_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][22] ),
    .C1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__a22o_1 _2202_ (.A1(\cpu.regFile.REGISTERS[10][22] ),
    .A2(_0459_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][22] ),
    .X(_0686_));
 sky130_fd_sc_hd__a211o_1 _2203_ (.A1(\cpu.regFile.REGISTERS[6][22] ),
    .A2(_0464_),
    .B1(_0686_),
    .C1(_0495_),
    .X(_0687_));
 sky130_fd_sc_hd__or3_2 _2204_ (.A(_0683_),
    .B(_0685_),
    .C(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__o221a_1 _2205_ (.A1(\cpu.regFile.REGISTERS[0][22] ),
    .A2(_0456_),
    .B1(_0681_),
    .B2(_0688_),
    .C1(_0499_),
    .X(_0689_));
 sky130_fd_sc_hd__a211o_1 _2206_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[22] ),
    .A2(_0454_),
    .B1(_0689_),
    .C1(_0502_),
    .X(_0690_));
 sky130_fd_sc_hd__o21ai_2 _2207_ (.A1(\cpu.ALU_OUT_MEMORY_4[22] ),
    .A2(_0450_),
    .B1(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__inv_2 _2208_ (.A(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__mux2_2 _2209_ (.A0(\cpu.immediateExtractor.VALUE[22] ),
    .A1(_0692_),
    .S(net126),
    .X(_0693_));
 sky130_fd_sc_hd__nor2_1 _2210_ (.A(_0679_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__mux2_1 _2211_ (.A0(\cpu.regFile.REGISTERS[0][21] ),
    .A1(\cpu.regFile.REGISTERS[6][21] ),
    .S(_0513_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _2212_ (.A0(net128),
    .A1(_0695_),
    .S(_0521_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(\cpu.ALU_OUT_MEMORY_4[21] ),
    .A1(_0696_),
    .S(_0527_),
    .X(_0697_));
 sky130_fd_sc_hd__and2_1 _2214_ (.A(_0509_),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__inv_2 _2215_ (.A(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__a22o_1 _2216_ (.A1(\cpu.regFile.REGISTERS[5][21] ),
    .A2(_0481_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][21] ),
    .X(_0700_));
 sky130_fd_sc_hd__a221o_1 _2217_ (.A1(\cpu.regFile.REGISTERS[11][21] ),
    .A2(_0461_),
    .B1(_0489_),
    .B2(\cpu.regFile.REGISTERS[12][21] ),
    .C1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__a22o_1 _2218_ (.A1(\cpu.regFile.REGISTERS[7][21] ),
    .A2(_0467_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][21] ),
    .X(_0702_));
 sky130_fd_sc_hd__a221o_1 _2219_ (.A1(\cpu.regFile.REGISTERS[15][21] ),
    .A2(_0469_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][21] ),
    .C1(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _2220_ (.A1(\cpu.regFile.REGISTERS[2][21] ),
    .A2(_0457_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][21] ),
    .X(_0704_));
 sky130_fd_sc_hd__a221o_1 _2221_ (.A1(\cpu.regFile.REGISTERS[3][21] ),
    .A2(_0471_),
    .B1(_0473_),
    .B2(\cpu.regFile.REGISTERS[14][21] ),
    .C1(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__a22o_1 _2222_ (.A1(\cpu.regFile.REGISTERS[10][21] ),
    .A2(_0459_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][21] ),
    .X(_0706_));
 sky130_fd_sc_hd__a211o_1 _2223_ (.A1(\cpu.regFile.REGISTERS[6][21] ),
    .A2(_0463_),
    .B1(_0706_),
    .C1(_0494_),
    .X(_0707_));
 sky130_fd_sc_hd__or3_2 _2224_ (.A(_0703_),
    .B(_0705_),
    .C(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__o221a_1 _2225_ (.A1(\cpu.regFile.REGISTERS[0][21] ),
    .A2(_0455_),
    .B1(_0701_),
    .B2(_0708_),
    .C1(_0498_),
    .X(_0709_));
 sky130_fd_sc_hd__a211o_1 _2226_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[21] ),
    .A2(_0453_),
    .B1(_0709_),
    .C1(_0501_),
    .X(_0710_));
 sky130_fd_sc_hd__o21a_1 _2227_ (.A1(\cpu.ALU_OUT_MEMORY_4[21] ),
    .A2(_0450_),
    .B1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _2228_ (.A0(\cpu.immediateExtractor.VALUE[21] ),
    .A1(_0711_),
    .S(net126),
    .X(_0712_));
 sky130_fd_sc_hd__nor2_1 _2229_ (.A(_0699_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(\cpu.regFile.REGISTERS[0][20] ),
    .A1(\cpu.regFile.REGISTERS[6][20] ),
    .S(_0513_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _2231_ (.A0(net117),
    .A1(_0714_),
    .S(_0521_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(\cpu.ALU_OUT_MEMORY_4[20] ),
    .A1(_0715_),
    .S(_0527_),
    .X(_0716_));
 sky130_fd_sc_hd__nand2_1 _2233_ (.A(_0509_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__a22o_1 _2234_ (.A1(\cpu.regFile.REGISTERS[5][20] ),
    .A2(_0481_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][20] ),
    .X(_0718_));
 sky130_fd_sc_hd__a221o_1 _2235_ (.A1(\cpu.regFile.REGISTERS[11][20] ),
    .A2(_0461_),
    .B1(_0489_),
    .B2(\cpu.regFile.REGISTERS[12][20] ),
    .C1(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__a22o_1 _2236_ (.A1(\cpu.regFile.REGISTERS[7][20] ),
    .A2(_0467_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][20] ),
    .X(_0720_));
 sky130_fd_sc_hd__a221o_1 _2237_ (.A1(\cpu.regFile.REGISTERS[15][20] ),
    .A2(_0469_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][20] ),
    .C1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__a22o_1 _2238_ (.A1(\cpu.regFile.REGISTERS[2][20] ),
    .A2(_0457_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][20] ),
    .X(_0722_));
 sky130_fd_sc_hd__a221o_1 _2239_ (.A1(\cpu.regFile.REGISTERS[3][20] ),
    .A2(_0471_),
    .B1(_0473_),
    .B2(\cpu.regFile.REGISTERS[14][20] ),
    .C1(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _2240_ (.A1(\cpu.regFile.REGISTERS[10][20] ),
    .A2(_0459_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][20] ),
    .X(_0724_));
 sky130_fd_sc_hd__a211o_1 _2241_ (.A1(\cpu.regFile.REGISTERS[6][20] ),
    .A2(_0463_),
    .B1(_0724_),
    .C1(_0494_),
    .X(_0725_));
 sky130_fd_sc_hd__or3_1 _2242_ (.A(_0721_),
    .B(_0723_),
    .C(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__o221a_1 _2243_ (.A1(\cpu.regFile.REGISTERS[0][20] ),
    .A2(_0455_),
    .B1(_0719_),
    .B2(_0726_),
    .C1(_0498_),
    .X(_0727_));
 sky130_fd_sc_hd__a211o_1 _2244_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[20] ),
    .A2(_0453_),
    .B1(_0727_),
    .C1(_0501_),
    .X(_0728_));
 sky130_fd_sc_hd__o21ai_2 _2245_ (.A1(\cpu.ALU_OUT_MEMORY_4[20] ),
    .A2(_0450_),
    .B1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_2 _2246_ (.A(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__mux2_2 _2247_ (.A0(\cpu.immediateExtractor.VALUE[20] ),
    .A1(_0730_),
    .S(net126),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _2248_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[19] ),
    .B(_0376_),
    .X(_0732_));
 sky130_fd_sc_hd__clkbuf_1 _2249_ (.A(_0732_),
    .X(\cpu.REG_WRITE_DATA[19] ));
 sky130_fd_sc_hd__mux2_1 _2250_ (.A0(\cpu.regFile.REGISTERS[0][19] ),
    .A1(\cpu.regFile.REGISTERS[6][19] ),
    .S(_0513_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _2251_ (.A0(net101),
    .A1(_0733_),
    .S(_0521_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _2252_ (.A0(\cpu.ALU_OUT_MEMORY_4[19] ),
    .A1(_0734_),
    .S(_0527_),
    .X(_0735_));
 sky130_fd_sc_hd__nand2_1 _2253_ (.A(_0509_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__inv_2 _2254_ (.A(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__a22o_1 _2255_ (.A1(\cpu.regFile.REGISTERS[11][19] ),
    .A2(_0461_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][19] ),
    .X(_0738_));
 sky130_fd_sc_hd__a221o_1 _2256_ (.A1(\cpu.regFile.REGISTERS[3][19] ),
    .A2(_0471_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][19] ),
    .C1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a22o_1 _2257_ (.A1(\cpu.regFile.REGISTERS[2][19] ),
    .A2(_0457_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][19] ),
    .X(_0740_));
 sky130_fd_sc_hd__a221o_1 _2258_ (.A1(\cpu.regFile.REGISTERS[5][19] ),
    .A2(_0481_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][19] ),
    .C1(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _2259_ (.A1(\cpu.regFile.REGISTERS[7][19] ),
    .A2(_0467_),
    .B1(_0459_),
    .B2(\cpu.regFile.REGISTERS[10][19] ),
    .X(_0742_));
 sky130_fd_sc_hd__a221o_1 _2260_ (.A1(\cpu.regFile.REGISTERS[12][19] ),
    .A2(_0489_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][19] ),
    .C1(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _2261_ (.A1(\cpu.regFile.REGISTERS[14][19] ),
    .A2(_0473_),
    .B1(_0469_),
    .B2(\cpu.regFile.REGISTERS[15][19] ),
    .X(_0744_));
 sky130_fd_sc_hd__a211o_1 _2262_ (.A1(\cpu.regFile.REGISTERS[6][19] ),
    .A2(_0463_),
    .B1(_0744_),
    .C1(_0494_),
    .X(_0745_));
 sky130_fd_sc_hd__or3_1 _2263_ (.A(_0741_),
    .B(_0743_),
    .C(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__o221a_1 _2264_ (.A1(\cpu.regFile.REGISTERS[0][19] ),
    .A2(_0455_),
    .B1(_0739_),
    .B2(_0746_),
    .C1(_0498_),
    .X(_0747_));
 sky130_fd_sc_hd__a211o_1 _2265_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[19] ),
    .A2(_0453_),
    .B1(_0747_),
    .C1(_0501_),
    .X(_0748_));
 sky130_fd_sc_hd__o21ai_4 _2266_ (.A1(\cpu.ALU_OUT_MEMORY_4[19] ),
    .A2(_0450_),
    .B1(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nor2_2 _2267_ (.A(_0536_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_1 _2268_ (.A(_0576_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__a2bb2o_1 _2269_ (.A1_N(_0717_),
    .A2_N(_0731_),
    .B1(_0737_),
    .B2(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__or3_1 _2270_ (.A(_0694_),
    .B(_0713_),
    .C(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _2271_ (.A1(\cpu.regFile.REGISTERS[1][16] ),
    .A2(_0487_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][16] ),
    .X(_0754_));
 sky130_fd_sc_hd__a221o_1 _2272_ (.A1(\cpu.regFile.REGISTERS[15][16] ),
    .A2(_0469_),
    .B1(_0489_),
    .B2(\cpu.regFile.REGISTERS[12][16] ),
    .C1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__a22o_1 _2273_ (.A1(\cpu.regFile.REGISTERS[11][16] ),
    .A2(_0461_),
    .B1(_0459_),
    .B2(\cpu.regFile.REGISTERS[10][16] ),
    .X(_0756_));
 sky130_fd_sc_hd__a221o_1 _2274_ (.A1(\cpu.regFile.REGISTERS[7][16] ),
    .A2(_0467_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][16] ),
    .C1(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__a22o_1 _2275_ (.A1(\cpu.regFile.REGISTERS[3][16] ),
    .A2(_0471_),
    .B1(_0481_),
    .B2(\cpu.regFile.REGISTERS[5][16] ),
    .X(_0758_));
 sky130_fd_sc_hd__a221o_1 _2276_ (.A1(\cpu.regFile.REGISTERS[2][16] ),
    .A2(_0457_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][16] ),
    .C1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__a22o_1 _2277_ (.A1(\cpu.regFile.REGISTERS[14][16] ),
    .A2(_0473_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][16] ),
    .X(_0760_));
 sky130_fd_sc_hd__a211o_1 _2278_ (.A1(\cpu.regFile.REGISTERS[6][16] ),
    .A2(_0463_),
    .B1(_0760_),
    .C1(_0494_),
    .X(_0761_));
 sky130_fd_sc_hd__or3_1 _2279_ (.A(_0757_),
    .B(_0759_),
    .C(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__o221a_1 _2280_ (.A1(\cpu.regFile.REGISTERS[0][16] ),
    .A2(_0455_),
    .B1(_0755_),
    .B2(_0762_),
    .C1(_0498_),
    .X(_0763_));
 sky130_fd_sc_hd__a211o_1 _2281_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[16] ),
    .A2(_0453_),
    .B1(_0763_),
    .C1(_0501_),
    .X(_0764_));
 sky130_fd_sc_hd__o21ai_4 _2282_ (.A1(\cpu.ALU_OUT_MEMORY_4[16] ),
    .A2(_0450_),
    .B1(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__nor2_1 _2283_ (.A(_0536_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__a21o_1 _2284_ (.A1(\cpu.immediateExtractor.VALUE[16] ),
    .A2(_0537_),
    .B1(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _2285_ (.A0(\cpu.regFile.REGISTERS[0][16] ),
    .A1(\cpu.regFile.REGISTERS[6][16] ),
    .S(_0513_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _2286_ (.A0(net113),
    .A1(_0768_),
    .S(_0521_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _2287_ (.A0(\cpu.ALU_OUT_MEMORY_4[16] ),
    .A1(_0769_),
    .S(_0527_),
    .X(_0770_));
 sky130_fd_sc_hd__nand2_1 _2288_ (.A(_0510_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__a22o_1 _2289_ (.A1(\cpu.regFile.REGISTERS[5][17] ),
    .A2(_0481_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][17] ),
    .X(_0772_));
 sky130_fd_sc_hd__a221o_1 _2290_ (.A1(\cpu.regFile.REGISTERS[12][17] ),
    .A2(_0489_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][17] ),
    .C1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _2291_ (.A1(\cpu.regFile.REGISTERS[11][17] ),
    .A2(_0240_),
    .B1(_0459_),
    .B2(\cpu.regFile.REGISTERS[10][17] ),
    .X(_0774_));
 sky130_fd_sc_hd__a221o_1 _2292_ (.A1(\cpu.regFile.REGISTERS[8][17] ),
    .A2(_0479_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][17] ),
    .C1(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__a22o_1 _2293_ (.A1(\cpu.regFile.REGISTERS[3][17] ),
    .A2(_0471_),
    .B1(_0469_),
    .B2(\cpu.regFile.REGISTERS[15][17] ),
    .X(_0776_));
 sky130_fd_sc_hd__a221o_1 _2294_ (.A1(\cpu.regFile.REGISTERS[2][17] ),
    .A2(_0457_),
    .B1(_0473_),
    .B2(\cpu.regFile.REGISTERS[14][17] ),
    .C1(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__a22o_1 _2295_ (.A1(\cpu.regFile.REGISTERS[7][17] ),
    .A2(_0301_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][17] ),
    .X(_0778_));
 sky130_fd_sc_hd__a211o_1 _2296_ (.A1(\cpu.regFile.REGISTERS[6][17] ),
    .A2(_0463_),
    .B1(_0778_),
    .C1(_0494_),
    .X(_0779_));
 sky130_fd_sc_hd__or3_1 _2297_ (.A(_0775_),
    .B(_0777_),
    .C(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o221a_1 _2298_ (.A1(\cpu.regFile.REGISTERS[0][17] ),
    .A2(_0455_),
    .B1(_0773_),
    .B2(_0780_),
    .C1(_0498_),
    .X(_0781_));
 sky130_fd_sc_hd__a211o_1 _2299_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[17] ),
    .A2(_0453_),
    .B1(_0781_),
    .C1(_0501_),
    .X(_0782_));
 sky130_fd_sc_hd__o21ai_1 _2300_ (.A1(\cpu.ALU_OUT_MEMORY_4[17] ),
    .A2(_0450_),
    .B1(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__inv_2 _2301_ (.A(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__mux2_1 _2302_ (.A0(\cpu.immediateExtractor.VALUE[16] ),
    .A1(_0784_),
    .S(net126),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _2303_ (.A0(\cpu.regFile.REGISTERS[0][17] ),
    .A1(\cpu.regFile.REGISTERS[6][17] ),
    .S(_0513_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _2304_ (.A0(net115),
    .A1(_0786_),
    .S(_0521_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _2305_ (.A0(\cpu.ALU_OUT_MEMORY_4[17] ),
    .A1(_0787_),
    .S(_0527_),
    .X(_0788_));
 sky130_fd_sc_hd__and2_1 _2306_ (.A(_0509_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__inv_2 _2307_ (.A(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__a22o_1 _2308_ (.A1(_0767_),
    .A2(_0771_),
    .B1(_0785_),
    .B2(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _2309_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[18] ),
    .B(_0376_),
    .X(_0792_));
 sky130_fd_sc_hd__clkbuf_1 _2310_ (.A(_0792_),
    .X(\cpu.REG_WRITE_DATA[18] ));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(\cpu.regFile.REGISTERS[0][18] ),
    .A1(\cpu.regFile.REGISTERS[6][18] ),
    .S(_0513_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _2312_ (.A0(net99),
    .A1(_0793_),
    .S(_0521_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _2313_ (.A0(\cpu.ALU_OUT_MEMORY_4[18] ),
    .A1(_0794_),
    .S(_0527_),
    .X(_0795_));
 sky130_fd_sc_hd__and2_2 _2314_ (.A(_0509_),
    .B(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__a22o_1 _2315_ (.A1(\cpu.regFile.REGISTERS[11][18] ),
    .A2(_0461_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][18] ),
    .X(_0797_));
 sky130_fd_sc_hd__a221o_1 _2316_ (.A1(\cpu.regFile.REGISTERS[3][18] ),
    .A2(_0472_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][18] ),
    .C1(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__a22o_1 _2317_ (.A1(\cpu.regFile.REGISTERS[2][18] ),
    .A2(_0457_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][18] ),
    .X(_0799_));
 sky130_fd_sc_hd__a221o_1 _2318_ (.A1(\cpu.regFile.REGISTERS[5][18] ),
    .A2(_0481_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][18] ),
    .C1(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_1 _2319_ (.A1(\cpu.regFile.REGISTERS[12][18] ),
    .A2(_0489_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][18] ),
    .X(_0801_));
 sky130_fd_sc_hd__a221o_1 _2320_ (.A1(\cpu.regFile.REGISTERS[7][18] ),
    .A2(_0468_),
    .B1(_0460_),
    .B2(\cpu.regFile.REGISTERS[10][18] ),
    .C1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _2321_ (.A1(\cpu.regFile.REGISTERS[14][18] ),
    .A2(_0473_),
    .B1(_0469_),
    .B2(\cpu.regFile.REGISTERS[15][18] ),
    .X(_0803_));
 sky130_fd_sc_hd__a211o_1 _2322_ (.A1(\cpu.regFile.REGISTERS[6][18] ),
    .A2(_0463_),
    .B1(_0803_),
    .C1(_0494_),
    .X(_0804_));
 sky130_fd_sc_hd__or3_1 _2323_ (.A(_0800_),
    .B(_0802_),
    .C(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__o221a_1 _2324_ (.A1(\cpu.regFile.REGISTERS[0][18] ),
    .A2(_0455_),
    .B1(_0798_),
    .B2(_0805_),
    .C1(_0498_),
    .X(_0806_));
 sky130_fd_sc_hd__a211o_1 _2325_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[18] ),
    .A2(_0453_),
    .B1(_0806_),
    .C1(_0501_),
    .X(_0807_));
 sky130_fd_sc_hd__o21ai_4 _2326_ (.A1(\cpu.ALU_OUT_MEMORY_4[18] ),
    .A2(_0450_),
    .B1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__o21a_2 _2327_ (.A1(_0536_),
    .A2(_0808_),
    .B1(_0551_),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _2328_ (.A(_0796_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nor2_1 _2329_ (.A(_0785_),
    .B(_0790_),
    .Y(_0811_));
 sky130_fd_sc_hd__or4_1 _2330_ (.A(_0753_),
    .B(_0791_),
    .C(_0810_),
    .D(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__a22o_1 _2331_ (.A1(_0699_),
    .A2(_0712_),
    .B1(_0717_),
    .B2(_0731_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _2332_ (.A0(\cpu.regFile.REGISTERS[0][23] ),
    .A1(\cpu.regFile.REGISTERS[6][23] ),
    .S(_0514_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(net121),
    .A1(_0814_),
    .S(_0522_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(\cpu.ALU_OUT_MEMORY_4[23] ),
    .A1(_0815_),
    .S(_0528_),
    .X(_0816_));
 sky130_fd_sc_hd__nand2_1 _2335_ (.A(_0510_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__a22o_1 _2336_ (.A1(\cpu.regFile.REGISTERS[5][23] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(\cpu.regFile.REGISTERS[13][23] ),
    .X(_0818_));
 sky130_fd_sc_hd__a221o_1 _2337_ (.A1(\cpu.regFile.REGISTERS[11][23] ),
    .A2(_0462_),
    .B1(_0490_),
    .B2(\cpu.regFile.REGISTERS[12][23] ),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _2338_ (.A1(\cpu.regFile.REGISTERS[7][23] ),
    .A2(_0468_),
    .B1(_0478_),
    .B2(\cpu.regFile.REGISTERS[9][23] ),
    .X(_0820_));
 sky130_fd_sc_hd__a221o_1 _2339_ (.A1(\cpu.regFile.REGISTERS[15][23] ),
    .A2(_0470_),
    .B1(_0480_),
    .B2(\cpu.regFile.REGISTERS[8][23] ),
    .C1(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__a22o_1 _2340_ (.A1(\cpu.regFile.REGISTERS[2][23] ),
    .A2(_0458_),
    .B1(_0488_),
    .B2(\cpu.regFile.REGISTERS[1][23] ),
    .X(_0822_));
 sky130_fd_sc_hd__a221o_1 _2341_ (.A1(\cpu.regFile.REGISTERS[3][23] ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(\cpu.regFile.REGISTERS[14][23] ),
    .C1(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__a22o_1 _2342_ (.A1(\cpu.regFile.REGISTERS[10][23] ),
    .A2(_0460_),
    .B1(_0492_),
    .B2(\cpu.regFile.REGISTERS[4][23] ),
    .X(_0824_));
 sky130_fd_sc_hd__a211o_1 _2343_ (.A1(\cpu.regFile.REGISTERS[6][23] ),
    .A2(_0464_),
    .B1(_0824_),
    .C1(_0495_),
    .X(_0825_));
 sky130_fd_sc_hd__or3_2 _2344_ (.A(_0821_),
    .B(_0823_),
    .C(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__o221a_1 _2345_ (.A1(\cpu.regFile.REGISTERS[0][23] ),
    .A2(_0456_),
    .B1(_0819_),
    .B2(_0826_),
    .C1(_0499_),
    .X(_0827_));
 sky130_fd_sc_hd__a211o_1 _2346_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[23] ),
    .A2(_0454_),
    .B1(_0827_),
    .C1(_0502_),
    .X(_0828_));
 sky130_fd_sc_hd__o21ai_4 _2347_ (.A1(\cpu.ALU_OUT_MEMORY_4[23] ),
    .A2(_0451_),
    .B1(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__o21ai_2 _2348_ (.A1(_0537_),
    .A2(_0829_),
    .B1(_0551_),
    .Y(_0830_));
 sky130_fd_sc_hd__a22o_1 _2349_ (.A1(_0679_),
    .A2(_0693_),
    .B1(_0817_),
    .B2(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__nor2_1 _2350_ (.A(_0737_),
    .B(_0751_),
    .Y(_0832_));
 sky130_fd_sc_hd__nor2_1 _2351_ (.A(_0817_),
    .B(_0830_),
    .Y(_0833_));
 sky130_fd_sc_hd__o22a_1 _2352_ (.A1(_0767_),
    .A2(_0771_),
    .B1(_0796_),
    .B2(_0809_),
    .X(_0834_));
 sky130_fd_sc_hd__or3b_1 _2353_ (.A(_0832_),
    .B(_0833_),
    .C_N(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__or4_1 _2354_ (.A(_0812_),
    .B(_0813_),
    .C(_0831_),
    .D(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _2355_ (.A(\cpu.REG_WRITE_DATA_WRITEBACK_5[14] ),
    .B(_0376_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _2356_ (.A(_0837_),
    .X(\cpu.REG_WRITE_DATA[14] ));
 sky130_fd_sc_hd__mux2_1 _2357_ (.A0(\cpu.regFile.REGISTERS[0][14] ),
    .A1(\cpu.regFile.REGISTERS[6][14] ),
    .S(_0513_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _2358_ (.A0(net97),
    .A1(_0838_),
    .S(_0521_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _2359_ (.A0(\cpu.ALU_OUT_MEMORY_4[14] ),
    .A1(_0839_),
    .S(_0527_),
    .X(_0840_));
 sky130_fd_sc_hd__and2_1 _2360_ (.A(_0509_),
    .B(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__a22o_1 _2361_ (.A1(\cpu.regFile.REGISTERS[11][14] ),
    .A2(_0461_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][14] ),
    .X(_0842_));
 sky130_fd_sc_hd__a221o_1 _2362_ (.A1(\cpu.regFile.REGISTERS[3][14] ),
    .A2(_0471_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][14] ),
    .C1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__a22o_1 _2363_ (.A1(\cpu.regFile.REGISTERS[5][14] ),
    .A2(_0481_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][14] ),
    .X(_0844_));
 sky130_fd_sc_hd__a221o_1 _2364_ (.A1(\cpu.regFile.REGISTERS[2][14] ),
    .A2(_0457_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][14] ),
    .C1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__a22o_1 _2365_ (.A1(\cpu.regFile.REGISTERS[7][14] ),
    .A2(_0467_),
    .B1(_0459_),
    .B2(\cpu.regFile.REGISTERS[10][14] ),
    .X(_0846_));
 sky130_fd_sc_hd__a221o_1 _2366_ (.A1(\cpu.regFile.REGISTERS[12][14] ),
    .A2(_0489_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][14] ),
    .C1(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__a22o_1 _2367_ (.A1(\cpu.regFile.REGISTERS[14][14] ),
    .A2(_0473_),
    .B1(_0469_),
    .B2(\cpu.regFile.REGISTERS[15][14] ),
    .X(_0848_));
 sky130_fd_sc_hd__a211o_1 _2368_ (.A1(\cpu.regFile.REGISTERS[6][14] ),
    .A2(_0463_),
    .B1(_0848_),
    .C1(_0494_),
    .X(_0849_));
 sky130_fd_sc_hd__or3_1 _2369_ (.A(_0845_),
    .B(_0847_),
    .C(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__o221a_1 _2370_ (.A1(\cpu.regFile.REGISTERS[0][14] ),
    .A2(_0455_),
    .B1(_0843_),
    .B2(_0850_),
    .C1(_0498_),
    .X(_0851_));
 sky130_fd_sc_hd__a211o_1 _2371_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[14] ),
    .A2(_0453_),
    .B1(_0851_),
    .C1(_0501_),
    .X(_0852_));
 sky130_fd_sc_hd__o21ai_4 _2372_ (.A1(\cpu.ALU_OUT_MEMORY_4[14] ),
    .A2(_0450_),
    .B1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__o21a_1 _2373_ (.A1(_0536_),
    .A2(_0853_),
    .B1(_0551_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(\cpu.regFile.REGISTERS[0][15] ),
    .A1(\cpu.regFile.REGISTERS[6][15] ),
    .S(_0513_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(net140),
    .A1(_0855_),
    .S(_0521_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(\cpu.ALU_OUT_MEMORY_4[15] ),
    .A1(_0856_),
    .S(_0527_),
    .X(_0857_));
 sky130_fd_sc_hd__nand2_1 _2377_ (.A(_0509_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a22o_1 _2378_ (.A1(\cpu.regFile.REGISTERS[10][15] ),
    .A2(_0459_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][15] ),
    .X(_0859_));
 sky130_fd_sc_hd__a221o_1 _2379_ (.A1(\cpu.regFile.REGISTERS[15][15] ),
    .A2(_0469_),
    .B1(_0463_),
    .B2(\cpu.regFile.REGISTERS[6][15] ),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a22o_1 _2380_ (.A1(\cpu.regFile.REGISTERS[3][15] ),
    .A2(_0471_),
    .B1(_0487_),
    .B2(\cpu.regFile.REGISTERS[1][15] ),
    .X(_0861_));
 sky130_fd_sc_hd__a221o_1 _2381_ (.A1(\cpu.regFile.REGISTERS[7][15] ),
    .A2(_0467_),
    .B1(_0489_),
    .B2(\cpu.regFile.REGISTERS[12][15] ),
    .C1(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__a22o_1 _2382_ (.A1(\cpu.regFile.REGISTERS[2][15] ),
    .A2(_0457_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][15] ),
    .X(_0863_));
 sky130_fd_sc_hd__a221o_1 _2383_ (.A1(\cpu.regFile.REGISTERS[11][15] ),
    .A2(_0461_),
    .B1(_0481_),
    .B2(\cpu.regFile.REGISTERS[5][15] ),
    .C1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__a22o_1 _2384_ (.A1(\cpu.regFile.REGISTERS[14][15] ),
    .A2(_0473_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][15] ),
    .X(_0865_));
 sky130_fd_sc_hd__a211o_1 _2385_ (.A1(\cpu.regFile.REGISTERS[8][15] ),
    .A2(_0479_),
    .B1(_0865_),
    .C1(_0494_),
    .X(_0866_));
 sky130_fd_sc_hd__or3_1 _2386_ (.A(_0862_),
    .B(_0864_),
    .C(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__o221a_1 _2387_ (.A1(\cpu.regFile.REGISTERS[0][15] ),
    .A2(_0455_),
    .B1(_0860_),
    .B2(_0867_),
    .C1(_0498_),
    .X(_0868_));
 sky130_fd_sc_hd__a211o_1 _2388_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[15] ),
    .A2(_0453_),
    .B1(_0868_),
    .C1(_0501_),
    .X(_0869_));
 sky130_fd_sc_hd__o21ai_4 _2389_ (.A1(\cpu.ALU_OUT_MEMORY_4[15] ),
    .A2(_0450_),
    .B1(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__o21ai_2 _2390_ (.A1(_0536_),
    .A2(_0870_),
    .B1(_0550_),
    .Y(_0871_));
 sky130_fd_sc_hd__a2bb2o_1 _2391_ (.A1_N(_0841_),
    .A2_N(_0854_),
    .B1(_0858_),
    .B2(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__inv_2 _2392_ (.A(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_1 _2393_ (.A(_0858_),
    .B(_0871_),
    .Y(_0874_));
 sky130_fd_sc_hd__mux2_1 _2394_ (.A0(\cpu.regFile.REGISTERS[0][13] ),
    .A1(\cpu.regFile.REGISTERS[6][13] ),
    .S(_0512_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(net138),
    .A1(_0875_),
    .S(_0520_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(\cpu.ALU_OUT_MEMORY_4[13] ),
    .A1(_0876_),
    .S(_0526_),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _2397_ (.A(_0510_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__a22o_1 _2398_ (.A1(\cpu.regFile.REGISTERS[10][13] ),
    .A2(_0459_),
    .B1(_0491_),
    .B2(\cpu.regFile.REGISTERS[4][13] ),
    .X(_0879_));
 sky130_fd_sc_hd__a221o_1 _2399_ (.A1(\cpu.regFile.REGISTERS[15][13] ),
    .A2(_0469_),
    .B1(_0463_),
    .B2(\cpu.regFile.REGISTERS[6][13] ),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__a22o_1 _2400_ (.A1(\cpu.regFile.REGISTERS[3][13] ),
    .A2(_0322_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][13] ),
    .X(_0881_));
 sky130_fd_sc_hd__a221o_1 _2401_ (.A1(\cpu.regFile.REGISTERS[7][13] ),
    .A2(_0467_),
    .B1(_0489_),
    .B2(\cpu.regFile.REGISTERS[12][13] ),
    .C1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _2402_ (.A1(\cpu.regFile.REGISTERS[2][13] ),
    .A2(_0305_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][13] ),
    .X(_0883_));
 sky130_fd_sc_hd__a221o_1 _2403_ (.A1(\cpu.regFile.REGISTERS[11][13] ),
    .A2(_0461_),
    .B1(_0481_),
    .B2(\cpu.regFile.REGISTERS[5][13] ),
    .C1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__a22o_1 _2404_ (.A1(\cpu.regFile.REGISTERS[14][13] ),
    .A2(_0291_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][13] ),
    .X(_0885_));
 sky130_fd_sc_hd__a211o_1 _2405_ (.A1(\cpu.regFile.REGISTERS[8][13] ),
    .A2(_0294_),
    .B1(_0885_),
    .C1(_0494_),
    .X(_0886_));
 sky130_fd_sc_hd__or3_2 _2406_ (.A(_0882_),
    .B(_0884_),
    .C(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__o221ai_4 _2407_ (.A1(\cpu.regFile.REGISTERS[0][13] ),
    .A2(_0455_),
    .B1(_0880_),
    .B2(_0887_),
    .C1(_0498_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21oi_1 _2408_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[13] ),
    .A2(_0452_),
    .B1(_0287_),
    .Y(_0889_));
 sky130_fd_sc_hd__a2bb2o_1 _2409_ (.A1_N(\cpu.ALU_OUT_MEMORY_4[13] ),
    .A2_N(_0342_),
    .B1(_0888_),
    .B2(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__clkinv_2 _2410_ (.A(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(\cpu.immediateExtractor.VALUE[13] ),
    .A1(_0891_),
    .S(_0012_),
    .X(_0892_));
 sky130_fd_sc_hd__a2bb2o_1 _2412_ (.A1_N(_0878_),
    .A2_N(_0892_),
    .B1(_0841_),
    .B2(_0854_),
    .X(_0893_));
 sky130_fd_sc_hd__or3_1 _2413_ (.A(_0872_),
    .B(_0874_),
    .C(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _2414_ (.A0(\cpu.regFile.REGISTERS[0][12] ),
    .A1(\cpu.regFile.REGISTERS[6][12] ),
    .S(_0513_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(net124),
    .A1(_0895_),
    .S(_0521_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_2 _2416_ (.A0(\cpu.ALU_OUT_MEMORY_4[12] ),
    .A1(_0896_),
    .S(_0527_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _2417_ (.A(_0510_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__a22o_1 _2418_ (.A1(\cpu.regFile.REGISTERS[14][12] ),
    .A2(_0473_),
    .B1(_0297_),
    .B2(\cpu.regFile.REGISTERS[4][12] ),
    .X(_0899_));
 sky130_fd_sc_hd__a221o_1 _2419_ (.A1(\cpu.regFile.REGISTERS[6][12] ),
    .A2(_0249_),
    .B1(_0479_),
    .B2(\cpu.regFile.REGISTERS[8][12] ),
    .C1(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__a22o_1 _2420_ (.A1(\cpu.regFile.REGISTERS[7][12] ),
    .A2(_0301_),
    .B1(_0314_),
    .B2(\cpu.regFile.REGISTERS[10][12] ),
    .X(_0901_));
 sky130_fd_sc_hd__a221o_1 _2421_ (.A1(\cpu.regFile.REGISTERS[3][12] ),
    .A2(_0322_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][12] ),
    .C1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_1 _2422_ (.A1(\cpu.regFile.REGISTERS[11][12] ),
    .A2(_0240_),
    .B1(_0305_),
    .B2(\cpu.regFile.REGISTERS[2][12] ),
    .X(_0903_));
 sky130_fd_sc_hd__a221o_1 _2423_ (.A1(\cpu.regFile.REGISTERS[15][12] ),
    .A2(_0247_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][12] ),
    .C1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _2424_ (.A1(\cpu.regFile.REGISTERS[9][12] ),
    .A2(_0292_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][12] ),
    .X(_0905_));
 sky130_fd_sc_hd__a211o_1 _2425_ (.A1(\cpu.regFile.REGISTERS[12][12] ),
    .A2(_0293_),
    .B1(_0905_),
    .C1(_0307_),
    .X(_0906_));
 sky130_fd_sc_hd__or3_2 _2426_ (.A(_0902_),
    .B(_0904_),
    .C(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__o221a_1 _2427_ (.A1(\cpu.regFile.REGISTERS[0][12] ),
    .A2(_0290_),
    .B1(_0900_),
    .B2(_0907_),
    .C1(_0289_),
    .X(_0908_));
 sky130_fd_sc_hd__a211o_1 _2428_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[12] ),
    .A2(_0453_),
    .B1(_0908_),
    .C1(_0501_),
    .X(_0909_));
 sky130_fd_sc_hd__o21ai_4 _2429_ (.A1(\cpu.ALU_OUT_MEMORY_4[12] ),
    .A2(_0342_),
    .B1(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__o21ai_2 _2430_ (.A1(_0536_),
    .A2(_0910_),
    .B1(_0550_),
    .Y(_0911_));
 sky130_fd_sc_hd__a22o_1 _2431_ (.A1(_0878_),
    .A2(_0892_),
    .B1(_0898_),
    .B2(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__inv_2 _2432_ (.A(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[7] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[7] ),
    .S(_0221_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2434_ (.A(_0914_),
    .X(\cpu.REG_WRITE_DATA[7] ));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(\cpu.regFile.REGISTERS[0][7] ),
    .A1(\cpu.regFile.REGISTERS[6][7] ),
    .S(_0512_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(net148),
    .A1(_0915_),
    .S(_0520_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_2 _2437_ (.A0(net177),
    .A1(_0916_),
    .S(_0526_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(\cpu.PC_EXECUTE_3[7] ),
    .A1(_0917_),
    .S(_0211_),
    .X(_0918_));
 sky130_fd_sc_hd__a22o_1 _2439_ (.A1(\cpu.regFile.REGISTERS[7][7] ),
    .A2(_0301_),
    .B1(_0314_),
    .B2(\cpu.regFile.REGISTERS[10][7] ),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _2440_ (.A1(\cpu.regFile.REGISTERS[15][7] ),
    .A2(_0247_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][7] ),
    .X(_0920_));
 sky130_fd_sc_hd__a22o_1 _2441_ (.A1(\cpu.regFile.REGISTERS[11][7] ),
    .A2(_0239_),
    .B1(_0248_),
    .B2(\cpu.regFile.REGISTERS[6][7] ),
    .X(_0921_));
 sky130_fd_sc_hd__a221o_1 _2442_ (.A1(\cpu.regFile.REGISTERS[3][7] ),
    .A2(_0322_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][7] ),
    .C1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__a22o_1 _2443_ (.A1(\cpu.regFile.REGISTERS[14][7] ),
    .A2(_0250_),
    .B1(_0264_),
    .B2(\cpu.regFile.REGISTERS[13][7] ),
    .X(_0923_));
 sky130_fd_sc_hd__a21o_1 _2444_ (.A1(\cpu.regFile.REGISTERS[1][7] ),
    .A2(_0302_),
    .B1(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _2445_ (.A1(\cpu.regFile.REGISTERS[12][7] ),
    .A2(_0254_),
    .B1(_0260_),
    .B2(\cpu.regFile.REGISTERS[4][7] ),
    .X(_0925_));
 sky130_fd_sc_hd__a21o_1 _2446_ (.A1(\cpu.regFile.REGISTERS[8][7] ),
    .A2(_0263_),
    .B1(_0261_),
    .X(_0926_));
 sky130_fd_sc_hd__a211o_1 _2447_ (.A1(\cpu.regFile.REGISTERS[2][7] ),
    .A2(_0305_),
    .B1(_0925_),
    .C1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__or4_2 _2448_ (.A(_0920_),
    .B(_0922_),
    .C(_0924_),
    .D(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__o221ai_2 _2449_ (.A1(\cpu.regFile.REGISTERS[0][7] ),
    .A2(_0290_),
    .B1(_0919_),
    .B2(_0928_),
    .C1(_0270_),
    .Y(_0929_));
 sky130_fd_sc_hd__a21oi_1 _2450_ (.A1(_0233_),
    .A2(net148),
    .B1(_0281_),
    .Y(_0930_));
 sky130_fd_sc_hd__a2bb2o_4 _2451_ (.A1_N(net176),
    .A2_N(_0342_),
    .B1(_0929_),
    .B2(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__or2_1 _2452_ (.A(_0506_),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__and2_1 _2453_ (.A(_0551_),
    .B(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _2454_ (.A0(\cpu.regFile.REGISTERS[0][8] ),
    .A1(\cpu.regFile.REGISTERS[6][8] ),
    .S(_0512_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(net130),
    .A1(_0934_),
    .S(_0520_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_2 _2456_ (.A0(net171),
    .A1(_0935_),
    .S(_0526_),
    .X(_0936_));
 sky130_fd_sc_hd__or2_1 _2457_ (.A(\cpu.PC_EXECUTE_3[8] ),
    .B(_0211_),
    .X(_0937_));
 sky130_fd_sc_hd__o21ai_2 _2458_ (.A1(_0206_),
    .A2(_0936_),
    .B1(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__a22o_1 _2459_ (.A1(\cpu.regFile.REGISTERS[14][8] ),
    .A2(_0291_),
    .B1(_0294_),
    .B2(\cpu.regFile.REGISTERS[8][8] ),
    .X(_0939_));
 sky130_fd_sc_hd__a221o_1 _2460_ (.A1(\cpu.regFile.REGISTERS[6][8] ),
    .A2(_0249_),
    .B1(_0483_),
    .B2(\cpu.regFile.REGISTERS[13][8] ),
    .C1(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__a22o_1 _2461_ (.A1(\cpu.regFile.REGISTERS[10][8] ),
    .A2(_0314_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][8] ),
    .X(_0941_));
 sky130_fd_sc_hd__a221o_1 _2462_ (.A1(\cpu.regFile.REGISTERS[2][8] ),
    .A2(_0457_),
    .B1(_0293_),
    .B2(\cpu.regFile.REGISTERS[12][8] ),
    .C1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__a22o_1 _2463_ (.A1(\cpu.regFile.REGISTERS[7][8] ),
    .A2(_0301_),
    .B1(_0297_),
    .B2(\cpu.regFile.REGISTERS[4][8] ),
    .X(_0943_));
 sky130_fd_sc_hd__a221o_1 _2464_ (.A1(\cpu.regFile.REGISTERS[15][8] ),
    .A2(_0247_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][8] ),
    .C1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__a22o_1 _2465_ (.A1(\cpu.regFile.REGISTERS[11][8] ),
    .A2(_0240_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][8] ),
    .X(_0945_));
 sky130_fd_sc_hd__a211o_1 _2466_ (.A1(\cpu.regFile.REGISTERS[3][8] ),
    .A2(_0471_),
    .B1(_0945_),
    .C1(_0307_),
    .X(_0946_));
 sky130_fd_sc_hd__or3_2 _2467_ (.A(_0942_),
    .B(_0944_),
    .C(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__o221ai_4 _2468_ (.A1(\cpu.regFile.REGISTERS[0][8] ),
    .A2(_0290_),
    .B1(_0940_),
    .B2(_0947_),
    .C1(_0289_),
    .Y(_0948_));
 sky130_fd_sc_hd__a21oi_1 _2469_ (.A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[8] ),
    .A2(_0452_),
    .B1(_0287_),
    .Y(_0949_));
 sky130_fd_sc_hd__a2bb2o_4 _2470_ (.A1_N(net170),
    .A2_N(_0342_),
    .B1(_0948_),
    .B2(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nor2_1 _2471_ (.A(_0536_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__or2_1 _2472_ (.A(_0576_),
    .B(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__o2bb2a_1 _2473_ (.A1_N(_0918_),
    .A2_N(_0933_),
    .B1(_0938_),
    .B2(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__clkinv_2 _2474_ (.A(\cpu.PC_EXECUTE_3[5] ),
    .Y(_0954_));
 sky130_fd_sc_hd__and4bb_2 _2475_ (.A_N(_0517_),
    .B_N(_0524_),
    .C(\cpu.R1_PIPELINE[1][1] ),
    .D(\cpu.RD_PIPELINE[2][1] ),
    .X(_0955_));
 sky130_fd_sc_hd__and4bb_1 _2476_ (.A_N(_0517_),
    .B_N(_0518_),
    .C(\cpu.R1_PIPELINE[1][1] ),
    .D(\cpu.RD_PIPELINE[3][1] ),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(\cpu.regFile.REGISTERS[0][5] ),
    .A1(\cpu.regFile.REGISTERS[6][5] ),
    .S(_0512_),
    .X(_0957_));
 sky130_fd_sc_hd__or2_1 _2478_ (.A(_0956_),
    .B(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__o211a_1 _2479_ (.A1(net143),
    .A2(_0520_),
    .B1(_0526_),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__a21oi_4 _2480_ (.A1(net188),
    .A2(_0955_),
    .B1(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__mux2_1 _2481_ (.A0(_0954_),
    .A1(_0960_),
    .S(_0510_),
    .X(_0961_));
 sky130_fd_sc_hd__a31o_1 _2482_ (.A1(_0346_),
    .A2(_0358_),
    .A3(_0507_),
    .B1(_0576_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(\cpu.regFile.REGISTERS[0][6] ),
    .A1(\cpu.regFile.REGISTERS[6][6] ),
    .S(\cpu.INSTRUCTION_EXECUTE_3[16] ),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _2484_ (.A(_0956_),
    .B(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__o211a_1 _2485_ (.A1(net152),
    .A2(_0519_),
    .B1(_0525_),
    .C1(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__a21oi_2 _2486_ (.A1(net183),
    .A2(_0955_),
    .B1(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__inv_2 _2487_ (.A(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(\cpu.PC_EXECUTE_3[6] ),
    .A1(_0967_),
    .S(_0211_),
    .X(_0968_));
 sky130_fd_sc_hd__a21oi_4 _2489_ (.A1(\cpu.R2_DATA[6] ),
    .A2(_0507_),
    .B1(_0576_),
    .Y(_0969_));
 sky130_fd_sc_hd__a2bb2o_1 _2490_ (.A1_N(_0961_),
    .A2_N(_0962_),
    .B1(_0968_),
    .B2(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_1 _2491_ (.A(\cpu.immediateExtractor.VALUE[4] ),
    .B(_0507_),
    .Y(_0971_));
 sky130_fd_sc_hd__a31o_1 _2492_ (.A1(_0361_),
    .A2(_0373_),
    .A3(_0507_),
    .B1(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_2 _2493_ (.A0(\cpu.regFile.REGISTERS[0][4] ),
    .A1(\cpu.regFile.REGISTERS[6][4] ),
    .S(_0512_),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(\cpu.REG_WRITE_DATA[4] ),
    .A1(_0973_),
    .S(_0520_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_2 _2495_ (.A0(net194),
    .A1(_0974_),
    .S(_0526_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(\cpu.PC_EXECUTE_3[4] ),
    .A1(_0975_),
    .S(_0211_),
    .X(_0976_));
 sky130_fd_sc_hd__and2_1 _2497_ (.A(_0972_),
    .B(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__nand2_1 _2498_ (.A(\cpu.immediateExtractor.VALUE[1] ),
    .B(_0506_),
    .Y(_0978_));
 sky130_fd_sc_hd__o31a_1 _2499_ (.A1(_0282_),
    .A2(_0284_),
    .A3(_0506_),
    .B1(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _2500_ (.A0(\cpu.regFile.REGISTERS[0][1] ),
    .A1(\cpu.regFile.REGISTERS[6][1] ),
    .S(\cpu.INSTRUCTION_EXECUTE_3[16] ),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(net160),
    .A1(_0980_),
    .S(_0519_),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(net212),
    .A1(_0981_),
    .S(_0525_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(\cpu.PC_EXECUTE_3[1] ),
    .A1(_0982_),
    .S(_0210_),
    .X(_0983_));
 sky130_fd_sc_hd__or2_1 _2504_ (.A(_0979_),
    .B(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__a22o_1 _2505_ (.A1(\cpu.regFile.REGISTERS[4][0] ),
    .A2(_0260_),
    .B1(_0264_),
    .B2(\cpu.regFile.REGISTERS[13][0] ),
    .X(_0985_));
 sky130_fd_sc_hd__a211o_1 _2506_ (.A1(\cpu.regFile.REGISTERS[3][0] ),
    .A2(_0322_),
    .B1(_0985_),
    .C1(_0307_),
    .X(_0986_));
 sky130_fd_sc_hd__a22o_1 _2507_ (.A1(\cpu.regFile.REGISTERS[11][0] ),
    .A2(_0239_),
    .B1(_0248_),
    .B2(\cpu.regFile.REGISTERS[6][0] ),
    .X(_0987_));
 sky130_fd_sc_hd__a221o_1 _2508_ (.A1(\cpu.regFile.REGISTERS[12][0] ),
    .A2(_0254_),
    .B1(_0263_),
    .B2(\cpu.regFile.REGISTERS[8][0] ),
    .C1(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__a22o_1 _2509_ (.A1(\cpu.regFile.REGISTERS[14][0] ),
    .A2(_0250_),
    .B1(_0246_),
    .B2(\cpu.regFile.REGISTERS[15][0] ),
    .X(_0989_));
 sky130_fd_sc_hd__a22o_1 _2510_ (.A1(\cpu.regFile.REGISTERS[10][0] ),
    .A2(_0251_),
    .B1(_0257_),
    .B2(\cpu.regFile.REGISTERS[9][0] ),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_1 _2511_ (.A1(\cpu.regFile.REGISTERS[7][0] ),
    .A2(_0238_),
    .B1(_0258_),
    .B2(\cpu.regFile.REGISTERS[5][0] ),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _2512_ (.A1(\cpu.regFile.REGISTERS[2][0] ),
    .A2(_0242_),
    .B1(_0255_),
    .B2(\cpu.regFile.REGISTERS[1][0] ),
    .X(_0992_));
 sky130_fd_sc_hd__or4_1 _2513_ (.A(_0989_),
    .B(_0990_),
    .C(_0991_),
    .D(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__or3_1 _2514_ (.A(_0986_),
    .B(_0988_),
    .C(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__or2_1 _2515_ (.A(\cpu.regFile.REGISTERS[0][0] ),
    .B(_0268_),
    .X(_0995_));
 sky130_fd_sc_hd__a21o_1 _2516_ (.A1(_0994_),
    .A2(_0995_),
    .B1(_0233_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(\cpu.RAM_READ_DATA_WRITEBACK_5[0] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[0] ),
    .S(_0221_),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(_0997_),
    .X(\cpu.REG_WRITE_DATA[0] ));
 sky130_fd_sc_hd__o21a_1 _2519_ (.A1(_0270_),
    .A2(net146),
    .B1(_0283_),
    .X(_0998_));
 sky130_fd_sc_hd__and2_1 _2520_ (.A(net218),
    .B(_0281_),
    .X(_0999_));
 sky130_fd_sc_hd__a21oi_4 _2521_ (.A1(_0996_),
    .A2(_0998_),
    .B1(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__nand2_1 _2522_ (.A(\cpu.immediateExtractor.VALUE[0] ),
    .B(_0506_),
    .Y(_1001_));
 sky130_fd_sc_hd__o21a_1 _2523_ (.A1(_0536_),
    .A2(_1000_),
    .B1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(\cpu.regFile.REGISTERS[0][0] ),
    .A1(\cpu.regFile.REGISTERS[6][0] ),
    .S(\cpu.INSTRUCTION_EXECUTE_3[16] ),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(net146),
    .A1(_1003_),
    .S(_0519_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(net219),
    .A1(_1004_),
    .S(_0525_),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(\cpu.PC_EXECUTE_3[0] ),
    .A1(_1005_),
    .S(_0210_),
    .X(_1006_));
 sky130_fd_sc_hd__nor2_1 _2528_ (.A(\cpu.immediateExtractor.VALUE[2] ),
    .B(_0507_),
    .Y(_1007_));
 sky130_fd_sc_hd__a31o_2 _2529_ (.A1(_0328_),
    .A2(_0329_),
    .A3(_0507_),
    .B1(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(\cpu.regFile.REGISTERS[0][2] ),
    .A1(\cpu.regFile.REGISTERS[6][2] ),
    .S(\cpu.INSTRUCTION_EXECUTE_3[16] ),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(net155),
    .A1(_1009_),
    .S(_0519_),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(net206),
    .A1(_1010_),
    .S(_0525_),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_2 _2533_ (.A0(\cpu.PC_EXECUTE_3[2] ),
    .A1(_1011_),
    .S(_0210_),
    .X(_1012_));
 sky130_fd_sc_hd__a22o_1 _2534_ (.A1(_1008_),
    .A2(_1012_),
    .B1(_0979_),
    .B2(_0983_),
    .X(_1013_));
 sky130_fd_sc_hd__nor2_1 _2535_ (.A(_1008_),
    .B(_1012_),
    .Y(_1014_));
 sky130_fd_sc_hd__nor2_1 _2536_ (.A(\cpu.immediateExtractor.VALUE[3] ),
    .B(_0507_),
    .Y(_1015_));
 sky130_fd_sc_hd__a31o_1 _2537_ (.A1(_0288_),
    .A2(_0312_),
    .A3(_0507_),
    .B1(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\cpu.regFile.REGISTERS[0][3] ),
    .A1(\cpu.regFile.REGISTERS[6][3] ),
    .S(_0512_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(\cpu.REG_WRITE_DATA[3] ),
    .A1(_1017_),
    .S(_0520_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_2 _2540_ (.A0(net200),
    .A1(_1018_),
    .S(_0526_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_2 _2541_ (.A0(\cpu.PC_EXECUTE_3[3] ),
    .A1(_1019_),
    .S(_0211_),
    .X(_1020_));
 sky130_fd_sc_hd__nor2_1 _2542_ (.A(_1016_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__nand2_1 _2543_ (.A(_1016_),
    .B(_1020_),
    .Y(_1022_));
 sky130_fd_sc_hd__or4b_1 _2544_ (.A(_1013_),
    .B(_1014_),
    .C(_1021_),
    .D_N(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__a31o_1 _2545_ (.A1(_0984_),
    .A2(_1002_),
    .A3(_1006_),
    .B1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__a21oi_1 _2546_ (.A1(_1014_),
    .A2(_1022_),
    .B1(_1021_),
    .Y(_1025_));
 sky130_fd_sc_hd__and2_1 _2547_ (.A(_1024_),
    .B(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__a2bb2o_1 _2548_ (.A1_N(_0972_),
    .A2_N(_0976_),
    .B1(_0962_),
    .B2(_0961_),
    .X(_1027_));
 sky130_fd_sc_hd__o21ba_1 _2549_ (.A1(_0977_),
    .A2(_1026_),
    .B1_N(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__o22a_1 _2550_ (.A1(_0933_),
    .A2(_0918_),
    .B1(_0969_),
    .B2(_0968_),
    .X(_1029_));
 sky130_fd_sc_hd__o21ai_1 _2551_ (.A1(_0970_),
    .A2(_1028_),
    .B1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(\cpu.regFile.REGISTERS[0][9] ),
    .A1(\cpu.regFile.REGISTERS[6][9] ),
    .S(_0512_),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(net132),
    .A1(_1031_),
    .S(_0520_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(net165),
    .A1(_1032_),
    .S(_0526_),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(\cpu.PC_EXECUTE_3[9] ),
    .A1(_1033_),
    .S(_0509_),
    .X(_1034_));
 sky130_fd_sc_hd__a22o_1 _2556_ (.A1(\cpu.regFile.REGISTERS[10][9] ),
    .A2(_0314_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][9] ),
    .X(_1035_));
 sky130_fd_sc_hd__a221o_1 _2557_ (.A1(\cpu.regFile.REGISTERS[7][9] ),
    .A2(_0467_),
    .B1(_0249_),
    .B2(\cpu.regFile.REGISTERS[6][9] ),
    .C1(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__a22o_1 _2558_ (.A1(\cpu.regFile.REGISTERS[2][9] ),
    .A2(_0305_),
    .B1(_0291_),
    .B2(\cpu.regFile.REGISTERS[14][9] ),
    .X(_1037_));
 sky130_fd_sc_hd__a221o_1 _2559_ (.A1(\cpu.regFile.REGISTERS[11][9] ),
    .A2(_0240_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][9] ),
    .C1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__a22o_1 _2560_ (.A1(\cpu.regFile.REGISTERS[15][9] ),
    .A2(_0247_),
    .B1(_0297_),
    .B2(\cpu.regFile.REGISTERS[4][9] ),
    .X(_1039_));
 sky130_fd_sc_hd__a211o_1 _2561_ (.A1(\cpu.regFile.REGISTERS[8][9] ),
    .A2(_0294_),
    .B1(_1039_),
    .C1(_0307_),
    .X(_1040_));
 sky130_fd_sc_hd__a22o_1 _2562_ (.A1(\cpu.regFile.REGISTERS[12][9] ),
    .A2(_0293_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][9] ),
    .X(_1041_));
 sky130_fd_sc_hd__a221o_1 _2563_ (.A1(\cpu.regFile.REGISTERS[3][9] ),
    .A2(_0322_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][9] ),
    .C1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__or3_2 _2564_ (.A(_1038_),
    .B(_1040_),
    .C(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__o21a_1 _2565_ (.A1(\cpu.regFile.REGISTERS[0][9] ),
    .A2(_0290_),
    .B1(_0289_),
    .X(_1044_));
 sky130_fd_sc_hd__o21ai_1 _2566_ (.A1(_1036_),
    .A2(_1043_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a21oi_1 _2567_ (.A1(_0233_),
    .A2(net132),
    .B1(_0287_),
    .Y(_1046_));
 sky130_fd_sc_hd__a2bb2o_2 _2568_ (.A1_N(net163),
    .A2_N(_0342_),
    .B1(_1045_),
    .B2(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__o21a_1 _2569_ (.A1(_0506_),
    .A2(_1047_),
    .B1(_0550_),
    .X(_1048_));
 sky130_fd_sc_hd__a2bb2o_1 _2570_ (.A1_N(_1034_),
    .A2_N(_1048_),
    .B1(_0938_),
    .B2(_0952_),
    .X(_1049_));
 sky130_fd_sc_hd__a21oi_1 _2571_ (.A1(_0953_),
    .A2(_1030_),
    .B1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(\cpu.regFile.REGISTERS[0][10] ),
    .A1(\cpu.regFile.REGISTERS[6][10] ),
    .S(_0512_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(\cpu.REG_WRITE_DATA[10] ),
    .A1(_1051_),
    .S(_0520_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_2 _2574_ (.A0(\cpu.ALU_OUT_MEMORY_4[10] ),
    .A1(_1052_),
    .S(_0526_),
    .X(_1053_));
 sky130_fd_sc_hd__and2_1 _2575_ (.A(_0511_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__a22o_1 _2576_ (.A1(\cpu.regFile.REGISTERS[12][10] ),
    .A2(_0293_),
    .B1(_0297_),
    .B2(\cpu.regFile.REGISTERS[4][10] ),
    .X(_1055_));
 sky130_fd_sc_hd__a221o_1 _2577_ (.A1(\cpu.regFile.REGISTERS[6][10] ),
    .A2(_0249_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][10] ),
    .C1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__a22o_1 _2578_ (.A1(\cpu.regFile.REGISTERS[3][10] ),
    .A2(_0322_),
    .B1(_0291_),
    .B2(\cpu.regFile.REGISTERS[14][10] ),
    .X(_1057_));
 sky130_fd_sc_hd__a221o_1 _2579_ (.A1(\cpu.regFile.REGISTERS[1][10] ),
    .A2(_0487_),
    .B1(_0477_),
    .B2(\cpu.regFile.REGISTERS[9][10] ),
    .C1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__a22o_1 _2580_ (.A1(\cpu.regFile.REGISTERS[7][10] ),
    .A2(_0301_),
    .B1(_0314_),
    .B2(\cpu.regFile.REGISTERS[10][10] ),
    .X(_1059_));
 sky130_fd_sc_hd__a22o_1 _2581_ (.A1(\cpu.regFile.REGISTERS[2][10] ),
    .A2(_0305_),
    .B1(_0247_),
    .B2(\cpu.regFile.REGISTERS[15][10] ),
    .X(_1060_));
 sky130_fd_sc_hd__a221o_1 _2582_ (.A1(\cpu.regFile.REGISTERS[11][10] ),
    .A2(_0240_),
    .B1(_0294_),
    .B2(\cpu.regFile.REGISTERS[8][10] ),
    .C1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__a2111o_1 _2583_ (.A1(\cpu.regFile.REGISTERS[13][10] ),
    .A2(_0298_),
    .B1(_1059_),
    .C1(_1061_),
    .D1(_0307_),
    .X(_1062_));
 sky130_fd_sc_hd__or3_1 _2584_ (.A(_1056_),
    .B(_1058_),
    .C(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__o211a_1 _2585_ (.A1(\cpu.regFile.REGISTERS[0][10] ),
    .A2(_0290_),
    .B1(_1063_),
    .C1(_0289_),
    .X(_1064_));
 sky130_fd_sc_hd__a21o_1 _2586_ (.A1(_0233_),
    .A2(\cpu.REG_WRITE_DATA[10] ),
    .B1(_0287_),
    .X(_1065_));
 sky130_fd_sc_hd__o22ai_4 _2587_ (.A1(\cpu.ALU_OUT_MEMORY_4[10] ),
    .A2(_0342_),
    .B1(_1064_),
    .B2(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__o21a_1 _2588_ (.A1(_0536_),
    .A2(_1066_),
    .B1(_0550_),
    .X(_1067_));
 sky130_fd_sc_hd__a22o_1 _2589_ (.A1(_1054_),
    .A2(_1067_),
    .B1(_1048_),
    .B2(_1034_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(\cpu.regFile.REGISTERS[0][11] ),
    .A1(\cpu.regFile.REGISTERS[6][11] ),
    .S(_0512_),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(\cpu.REG_WRITE_DATA[11] ),
    .A1(_1069_),
    .S(_0520_),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(\cpu.ALU_OUT_MEMORY_4[11] ),
    .A1(_1070_),
    .S(_0526_),
    .X(_1071_));
 sky130_fd_sc_hd__and2_1 _2593_ (.A(_0211_),
    .B(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__clkinv_2 _2594_ (.A(\cpu.immediateExtractor.VALUE[11] ),
    .Y(_1073_));
 sky130_fd_sc_hd__a22o_1 _2595_ (.A1(\cpu.regFile.REGISTERS[2][11] ),
    .A2(_0305_),
    .B1(_0291_),
    .B2(\cpu.regFile.REGISTERS[14][11] ),
    .X(_1074_));
 sky130_fd_sc_hd__a221o_1 _2596_ (.A1(\cpu.regFile.REGISTERS[11][11] ),
    .A2(_0461_),
    .B1(_0292_),
    .B2(\cpu.regFile.REGISTERS[9][11] ),
    .C1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__a22o_1 _2597_ (.A1(\cpu.regFile.REGISTERS[10][11] ),
    .A2(_0314_),
    .B1(_0298_),
    .B2(\cpu.regFile.REGISTERS[13][11] ),
    .X(_1076_));
 sky130_fd_sc_hd__a221o_1 _2598_ (.A1(\cpu.regFile.REGISTERS[7][11] ),
    .A2(_0301_),
    .B1(_0249_),
    .B2(\cpu.regFile.REGISTERS[6][11] ),
    .C1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__a22o_1 _2599_ (.A1(\cpu.regFile.REGISTERS[15][11] ),
    .A2(_0247_),
    .B1(_0297_),
    .B2(\cpu.regFile.REGISTERS[4][11] ),
    .X(_1078_));
 sky130_fd_sc_hd__a22o_1 _2600_ (.A1(\cpu.regFile.REGISTERS[3][11] ),
    .A2(_0322_),
    .B1(_0317_),
    .B2(\cpu.regFile.REGISTERS[5][11] ),
    .X(_1079_));
 sky130_fd_sc_hd__a221o_1 _2601_ (.A1(\cpu.regFile.REGISTERS[12][11] ),
    .A2(_0293_),
    .B1(_0302_),
    .B2(\cpu.regFile.REGISTERS[1][11] ),
    .C1(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__a2111o_1 _2602_ (.A1(\cpu.regFile.REGISTERS[8][11] ),
    .A2(_0294_),
    .B1(_1078_),
    .C1(_1080_),
    .D1(_0307_),
    .X(_1081_));
 sky130_fd_sc_hd__or3_1 _2603_ (.A(_1075_),
    .B(_1077_),
    .C(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__o211ai_2 _2604_ (.A1(\cpu.regFile.REGISTERS[0][11] ),
    .A2(_0290_),
    .B1(_1082_),
    .C1(_0289_),
    .Y(_1083_));
 sky130_fd_sc_hd__a21oi_1 _2605_ (.A1(_0233_),
    .A2(\cpu.REG_WRITE_DATA[11] ),
    .B1(_0287_),
    .Y(_1084_));
 sky130_fd_sc_hd__a2bb2o_2 _2606_ (.A1_N(\cpu.ALU_OUT_MEMORY_4[11] ),
    .A2_N(_0342_),
    .B1(_1083_),
    .B2(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(_1073_),
    .A1(_1085_),
    .S(net125),
    .X(_1086_));
 sky130_fd_sc_hd__o22a_1 _2608_ (.A1(_1054_),
    .A2(_1067_),
    .B1(_1072_),
    .B2(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__o21a_1 _2609_ (.A1(_1050_),
    .A2(_1068_),
    .B1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__inv_2 _2610_ (.A(_0911_),
    .Y(_1089_));
 sky130_fd_sc_hd__a311o_1 _2611_ (.A1(_0511_),
    .A2(_0897_),
    .A3(_1089_),
    .B1(_0912_),
    .C1(_0894_),
    .X(_1090_));
 sky130_fd_sc_hd__and2_1 _2612_ (.A(_1072_),
    .B(_1086_),
    .X(_1091_));
 sky130_fd_sc_hd__or3_1 _2613_ (.A(_1088_),
    .B(_1090_),
    .C(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__o221a_1 _2614_ (.A1(_0873_),
    .A2(_0874_),
    .B1(_0894_),
    .B2(_0913_),
    .C1(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__clkinv_2 _2615_ (.A(_0791_),
    .Y(_1094_));
 sky130_fd_sc_hd__or3_1 _2616_ (.A(_1094_),
    .B(_0810_),
    .C(_0811_),
    .X(_1095_));
 sky130_fd_sc_hd__o221a_1 _2617_ (.A1(_0737_),
    .A2(_0751_),
    .B1(_0796_),
    .B2(_0809_),
    .C1(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__o21ba_1 _2618_ (.A1(_0752_),
    .A2(_1096_),
    .B1_N(_0813_),
    .X(_1097_));
 sky130_fd_sc_hd__inv_2 _2619_ (.A(_0831_),
    .Y(_1098_));
 sky130_fd_sc_hd__o31a_1 _2620_ (.A1(_0694_),
    .A2(_0713_),
    .A3(_1097_),
    .B1(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__o22a_1 _2621_ (.A1(_0836_),
    .A2(_1093_),
    .B1(_1099_),
    .B2(_0833_),
    .X(_1100_));
 sky130_fd_sc_hd__o22a_1 _2622_ (.A1(_0592_),
    .A2(_0594_),
    .B1(_0595_),
    .B2(_0653_),
    .X(_1101_));
 sky130_fd_sc_hd__o21ba_1 _2623_ (.A1(_0633_),
    .A2(_1101_),
    .B1_N(_0632_),
    .X(_1102_));
 sky130_fd_sc_hd__o21ba_1 _2624_ (.A1(_0674_),
    .A2(_1102_),
    .B1_N(_0673_),
    .X(_1103_));
 sky130_fd_sc_hd__o21ai_1 _2625_ (.A1(_0675_),
    .A2(_1100_),
    .B1(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__and4bb_1 _2626_ (.A_N(_1049_),
    .B_N(_0977_),
    .C(_0984_),
    .D(_1029_),
    .X(_1105_));
 sky130_fd_sc_hd__nand2_1 _2627_ (.A(_0953_),
    .B(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__or3_1 _2628_ (.A(_0836_),
    .B(_1090_),
    .C(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__nand2_1 _2629_ (.A(_1002_),
    .B(_1006_),
    .Y(_1108_));
 sky130_fd_sc_hd__or2_1 _2630_ (.A(_1002_),
    .B(_1006_),
    .X(_1109_));
 sky130_fd_sc_hd__nand2_1 _2631_ (.A(_1108_),
    .B(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__or4b_1 _2632_ (.A(_1023_),
    .B(_1091_),
    .C(_1068_),
    .D_N(_1087_),
    .X(_1111_));
 sky130_fd_sc_hd__or4_1 _2633_ (.A(_0970_),
    .B(_1027_),
    .C(_1110_),
    .D(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_4 _2634_ (.A(_0207_),
    .X(_1113_));
 sky130_fd_sc_hd__and4b_1 _2635_ (.A_N(_1113_),
    .B(\cpu.INSTRUCTION_EXECUTE_3[13] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[0] ),
    .D(\cpu.INSTRUCTION_EXECUTE_3[4] ),
    .X(_1114_));
 sky130_fd_sc_hd__buf_4 _2636_ (.A(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__o31a_1 _2637_ (.A1(_0675_),
    .A2(_1107_),
    .A3(_1112_),
    .B1(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__nand4b_4 _2638_ (.A_N(_1113_),
    .B(\cpu.INSTRUCTION_EXECUTE_3[13] ),
    .C(\cpu.INSTRUCTION_EXECUTE_3[0] ),
    .D(\cpu.INSTRUCTION_EXECUTE_3[4] ),
    .Y(_1117_));
 sky130_fd_sc_hd__clkbuf_8 _2639_ (.A(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__a32o_1 _2640_ (.A1(_0531_),
    .A2(_1104_),
    .A3(_1116_),
    .B1(_1118_),
    .B2(_1110_),
    .X(_0163_));
 sky130_fd_sc_hd__o211a_2 _2641_ (.A1(_0506_),
    .A2(_1000_),
    .B1(_1001_),
    .C1(_0979_),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_1 _2642_ (.A(\cpu.immediateExtractor.VALUE[0] ),
    .B(net125),
    .Y(_1120_));
 sky130_fd_sc_hd__a211oi_1 _2643_ (.A1(net125),
    .A2(_1000_),
    .B1(_1120_),
    .C1(_0979_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21a_1 _2644_ (.A1(_1119_),
    .A2(_1121_),
    .B1(_0983_),
    .X(_1122_));
 sky130_fd_sc_hd__or3_1 _2645_ (.A(_0983_),
    .B(_1119_),
    .C(_1121_),
    .X(_1123_));
 sky130_fd_sc_hd__and2b_1 _2646_ (.A_N(_1122_),
    .B(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__buf_6 _2647_ (.A(_1115_),
    .X(_1125_));
 sky130_fd_sc_hd__a21oi_1 _2648_ (.A1(_1109_),
    .A2(_1124_),
    .B1(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__o21a_1 _2649_ (.A1(_1109_),
    .A2(_1124_),
    .B1(_1126_),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_1 _2650_ (.A1(_1109_),
    .A2(_1123_),
    .B1(_1122_),
    .X(_1127_));
 sky130_fd_sc_hd__xnor2_1 _2651_ (.A(_1008_),
    .B(_1119_),
    .Y(_1128_));
 sky130_fd_sc_hd__xor2_2 _2652_ (.A(_1012_),
    .B(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__a21oi_1 _2653_ (.A1(_1127_),
    .A2(_1129_),
    .B1(_1125_),
    .Y(_1130_));
 sky130_fd_sc_hd__o21a_1 _2654_ (.A1(_1127_),
    .A2(_1129_),
    .B1(_1130_),
    .X(_0185_));
 sky130_fd_sc_hd__and3_1 _2655_ (.A(_1008_),
    .B(_1016_),
    .C(_1119_),
    .X(_1131_));
 sky130_fd_sc_hd__a21oi_1 _2656_ (.A1(_1008_),
    .A2(_1119_),
    .B1(_1016_),
    .Y(_1132_));
 sky130_fd_sc_hd__or2_1 _2657_ (.A(_1131_),
    .B(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__or2_1 _2658_ (.A(_1020_),
    .B(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _2659_ (.A(_1020_),
    .B(_1133_),
    .Y(_1135_));
 sky130_fd_sc_hd__and2_1 _2660_ (.A(_1012_),
    .B(_1128_),
    .X(_1136_));
 sky130_fd_sc_hd__a21o_1 _2661_ (.A1(_1127_),
    .A2(_1129_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__a21oi_1 _2662_ (.A1(_1134_),
    .A2(_1135_),
    .B1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__a31o_1 _2663_ (.A1(_1134_),
    .A2(_1135_),
    .A3(_1137_),
    .B1(_1115_),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_1 _2664_ (.A(_1138_),
    .B(_1139_),
    .Y(_0188_));
 sky130_fd_sc_hd__xnor2_1 _2665_ (.A(_0972_),
    .B(_1131_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _2666_ (.A(_0976_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__or2_1 _2667_ (.A(_0976_),
    .B(_1140_),
    .X(_1142_));
 sky130_fd_sc_hd__and2_1 _2668_ (.A(_1141_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nor2_1 _2669_ (.A(_1020_),
    .B(_1133_),
    .Y(_1144_));
 sky130_fd_sc_hd__a221oi_2 _2670_ (.A1(_1127_),
    .A2(_1129_),
    .B1(_1133_),
    .B2(_1020_),
    .C1(_1136_),
    .Y(_1145_));
 sky130_fd_sc_hd__nor2_1 _2671_ (.A(_1144_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__a21oi_1 _2672_ (.A1(_1143_),
    .A2(_1146_),
    .B1(_1125_),
    .Y(_1147_));
 sky130_fd_sc_hd__o21a_1 _2673_ (.A1(_1143_),
    .A2(_1146_),
    .B1(_1147_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _2674_ (.A(_0960_),
    .Y(_1148_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(\cpu.PC_EXECUTE_3[5] ),
    .A1(_1148_),
    .S(_0211_),
    .X(_1149_));
 sky130_fd_sc_hd__and4_1 _2676_ (.A(_0972_),
    .B(_1008_),
    .C(_1016_),
    .D(_1119_),
    .X(_1150_));
 sky130_fd_sc_hd__xor2_1 _2677_ (.A(_0962_),
    .B(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__and2_1 _2678_ (.A(_1149_),
    .B(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__nor2_1 _2679_ (.A(_1149_),
    .B(_1151_),
    .Y(_1153_));
 sky130_fd_sc_hd__nor2_1 _2680_ (.A(_1152_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a21bo_1 _2681_ (.A1(_1143_),
    .A2(_1146_),
    .B1_N(_1141_),
    .X(_1155_));
 sky130_fd_sc_hd__nand2_1 _2682_ (.A(_1154_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__o211a_1 _2683_ (.A1(_1154_),
    .A2(_1155_),
    .B1(_1156_),
    .C1(_1118_),
    .X(_0190_));
 sky130_fd_sc_hd__and2b_1 _2684_ (.A_N(_0962_),
    .B(_0972_),
    .X(_1157_));
 sky130_fd_sc_hd__a21oi_1 _2685_ (.A1(_1131_),
    .A2(_1157_),
    .B1(_0969_),
    .Y(_1158_));
 sky130_fd_sc_hd__and3_1 _2686_ (.A(_0969_),
    .B(_1131_),
    .C(_1157_),
    .X(_1159_));
 sky130_fd_sc_hd__o21a_1 _2687_ (.A1(_1158_),
    .A2(_1159_),
    .B1(_0968_),
    .X(_1160_));
 sky130_fd_sc_hd__or3_1 _2688_ (.A(_0968_),
    .B(_1158_),
    .C(_1159_),
    .X(_1161_));
 sky130_fd_sc_hd__or2b_1 _2689_ (.A(_1160_),
    .B_N(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__xnor2_1 _2690_ (.A(_0976_),
    .B(_1140_),
    .Y(_1163_));
 sky130_fd_sc_hd__nand2_1 _2691_ (.A(_1149_),
    .B(_1151_),
    .Y(_1164_));
 sky130_fd_sc_hd__o311a_1 _2692_ (.A1(_1144_),
    .A2(_1163_),
    .A3(_1145_),
    .B1(_1164_),
    .C1(_1141_),
    .X(_1165_));
 sky130_fd_sc_hd__or2_1 _2693_ (.A(_1153_),
    .B(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__o21ai_1 _2694_ (.A1(_1162_),
    .A2(_1166_),
    .B1(_1118_),
    .Y(_1167_));
 sky130_fd_sc_hd__a21oi_1 _2695_ (.A1(_1162_),
    .A2(_1166_),
    .B1(_1167_),
    .Y(_0191_));
 sky130_fd_sc_hd__and4_1 _2696_ (.A(_0932_),
    .B(_1008_),
    .C(_1016_),
    .D(_1119_),
    .X(_1168_));
 sky130_fd_sc_hd__and3_1 _2697_ (.A(_0969_),
    .B(_1157_),
    .C(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__buf_2 _2698_ (.A(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__a31oi_1 _2699_ (.A1(_0969_),
    .A2(_1131_),
    .A3(_1157_),
    .B1(_0933_),
    .Y(_1171_));
 sky130_fd_sc_hd__or3_1 _2700_ (.A(_0918_),
    .B(_1170_),
    .C(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__o21ai_1 _2701_ (.A1(_1170_),
    .A2(_1171_),
    .B1(_0918_),
    .Y(_1173_));
 sky130_fd_sc_hd__nand2_1 _2702_ (.A(_1172_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__o21ba_1 _2703_ (.A1(_1162_),
    .A2(_1166_),
    .B1_N(_1160_),
    .X(_1175_));
 sky130_fd_sc_hd__nor2_1 _2704_ (.A(_1174_),
    .B(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__a211oi_1 _2705_ (.A1(_1174_),
    .A2(_1175_),
    .B1(_1176_),
    .C1(_1125_),
    .Y(_0192_));
 sky130_fd_sc_hd__xnor2_1 _2706_ (.A(_0952_),
    .B(_1170_),
    .Y(_1177_));
 sky130_fd_sc_hd__xor2_1 _2707_ (.A(_0938_),
    .B(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__inv_2 _2708_ (.A(_1172_),
    .Y(_1179_));
 sky130_fd_sc_hd__and2b_1 _2709_ (.A_N(_1160_),
    .B(_1173_),
    .X(_1180_));
 sky130_fd_sc_hd__o31a_1 _2710_ (.A1(_1153_),
    .A2(_1162_),
    .A3(_1165_),
    .B1(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__nor2_1 _2711_ (.A(_1179_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__and2_1 _2712_ (.A(_1178_),
    .B(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__o21ai_1 _2713_ (.A1(_1178_),
    .A2(_1182_),
    .B1(_1118_),
    .Y(_1184_));
 sky130_fd_sc_hd__nor2_1 _2714_ (.A(_1183_),
    .B(_1184_),
    .Y(_0193_));
 sky130_fd_sc_hd__nor2_1 _2715_ (.A(_0938_),
    .B(_1177_),
    .Y(_1185_));
 sky130_fd_sc_hd__and2b_1 _2716_ (.A_N(_0951_),
    .B(_1048_),
    .X(_1186_));
 sky130_fd_sc_hd__nor2_1 _2717_ (.A(_0576_),
    .B(_0951_),
    .Y(_1187_));
 sky130_fd_sc_hd__a41o_1 _2718_ (.A1(_1187_),
    .A2(_0969_),
    .A3(_1157_),
    .A4(_1168_),
    .B1(_1048_),
    .X(_1188_));
 sky130_fd_sc_hd__a21bo_1 _2719_ (.A1(_1170_),
    .A2(_1186_),
    .B1_N(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__xor2_1 _2720_ (.A(_1034_),
    .B(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__o21ai_1 _2721_ (.A1(_1185_),
    .A2(_1183_),
    .B1(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__or3_1 _2722_ (.A(_1185_),
    .B(_1183_),
    .C(_1190_),
    .X(_1192_));
 sky130_fd_sc_hd__and3_1 _2723_ (.A(_1117_),
    .B(_1191_),
    .C(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2724_ (.A(_1193_),
    .X(_0194_));
 sky130_fd_sc_hd__nand3_1 _2725_ (.A(_1067_),
    .B(_1170_),
    .C(_1186_),
    .Y(_1194_));
 sky130_fd_sc_hd__a21o_1 _2726_ (.A1(_1170_),
    .A2(_1186_),
    .B1(_1067_),
    .X(_1195_));
 sky130_fd_sc_hd__nand2_1 _2727_ (.A(_0211_),
    .B(_1053_),
    .Y(_1196_));
 sky130_fd_sc_hd__a21oi_2 _2728_ (.A1(_1194_),
    .A2(_1195_),
    .B1(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__and3_1 _2729_ (.A(_1196_),
    .B(_1194_),
    .C(_1195_),
    .X(_1198_));
 sky130_fd_sc_hd__nor2_2 _2730_ (.A(_1197_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__a21o_1 _2731_ (.A1(_1034_),
    .A2(_1189_),
    .B1(_1185_),
    .X(_1200_));
 sky130_fd_sc_hd__or2_1 _2732_ (.A(_1034_),
    .B(_1189_),
    .X(_1201_));
 sky130_fd_sc_hd__o21a_1 _2733_ (.A1(_1183_),
    .A2(_1200_),
    .B1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__o21ai_1 _2734_ (.A1(_1199_),
    .A2(_1202_),
    .B1(_1118_),
    .Y(_1203_));
 sky130_fd_sc_hd__a21oi_1 _2735_ (.A1(_1199_),
    .A2(_1202_),
    .B1(_1203_),
    .Y(_0164_));
 sky130_fd_sc_hd__and3_1 _2736_ (.A(_1067_),
    .B(_1086_),
    .C(_1186_),
    .X(_1204_));
 sky130_fd_sc_hd__and2_1 _2737_ (.A(_1170_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__a31oi_1 _2738_ (.A1(_1067_),
    .A2(_1170_),
    .A3(_1186_),
    .B1(_1086_),
    .Y(_1206_));
 sky130_fd_sc_hd__nor3_1 _2739_ (.A(_1072_),
    .B(_1205_),
    .C(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__o21a_1 _2740_ (.A1(_1205_),
    .A2(_1206_),
    .B1(_1072_),
    .X(_1208_));
 sky130_fd_sc_hd__or2_1 _2741_ (.A(_1207_),
    .B(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__a21oi_1 _2742_ (.A1(_1199_),
    .A2(_1202_),
    .B1(_1197_),
    .Y(_1210_));
 sky130_fd_sc_hd__a21oi_1 _2743_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1125_),
    .Y(_1211_));
 sky130_fd_sc_hd__o21a_1 _2744_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1211_),
    .X(_0165_));
 sky130_fd_sc_hd__or4_1 _2745_ (.A(_1197_),
    .B(_1198_),
    .C(_1207_),
    .D(_1208_),
    .X(_1212_));
 sky130_fd_sc_hd__nand2_1 _2746_ (.A(_1178_),
    .B(_1190_),
    .Y(_1213_));
 sky130_fd_sc_hd__or4_2 _2747_ (.A(_1179_),
    .B(_1181_),
    .C(_1212_),
    .D(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_1 _2748_ (.A(_1207_),
    .B(_1208_),
    .Y(_1215_));
 sky130_fd_sc_hd__o21ba_1 _2749_ (.A1(_1197_),
    .A2(_1208_),
    .B1_N(_1207_),
    .X(_1216_));
 sky130_fd_sc_hd__a41oi_4 _2750_ (.A1(_1201_),
    .A2(_1199_),
    .A3(_1200_),
    .A4(_1215_),
    .B1(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__xnor2_2 _2751_ (.A(_0911_),
    .B(_1205_),
    .Y(_1218_));
 sky130_fd_sc_hd__xnor2_1 _2752_ (.A(_0898_),
    .B(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__a21oi_1 _2753_ (.A1(_1214_),
    .A2(_1217_),
    .B1(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a31o_1 _2754_ (.A1(_1219_),
    .A2(_1214_),
    .A3(_1217_),
    .B1(_1115_),
    .X(_1221_));
 sky130_fd_sc_hd__nor2_1 _2755_ (.A(_1220_),
    .B(_1221_),
    .Y(_0166_));
 sky130_fd_sc_hd__and4b_1 _2756_ (.A_N(_0892_),
    .B(_1089_),
    .C(_1170_),
    .D(_1204_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_2 _2757_ (.A(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__a21boi_1 _2758_ (.A1(_1089_),
    .A2(_1205_),
    .B1_N(_0892_),
    .Y(_1224_));
 sky130_fd_sc_hd__and2_1 _2759_ (.A(_0509_),
    .B(_0877_),
    .X(_1225_));
 sky130_fd_sc_hd__o21ai_1 _2760_ (.A1(_1223_),
    .A2(_1224_),
    .B1(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__or3_1 _2761_ (.A(_1225_),
    .B(_1223_),
    .C(_1224_),
    .X(_1227_));
 sky130_fd_sc_hd__nand2_1 _2762_ (.A(_1226_),
    .B(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__o21ba_1 _2763_ (.A1(_0898_),
    .A2(_1218_),
    .B1_N(_1220_),
    .X(_1229_));
 sky130_fd_sc_hd__a21oi_1 _2764_ (.A1(_1228_),
    .A2(_1229_),
    .B1(_1125_),
    .Y(_1230_));
 sky130_fd_sc_hd__o21a_1 _2765_ (.A1(_1228_),
    .A2(_1229_),
    .B1(_1230_),
    .X(_0167_));
 sky130_fd_sc_hd__o21ai_1 _2766_ (.A1(_0898_),
    .A2(_1218_),
    .B1(_1226_),
    .Y(_1231_));
 sky130_fd_sc_hd__or2_1 _2767_ (.A(_1220_),
    .B(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__o21ai_1 _2768_ (.A1(_0537_),
    .A2(_0853_),
    .B1(_0551_),
    .Y(_1233_));
 sky130_fd_sc_hd__xnor2_1 _2769_ (.A(_1233_),
    .B(_1223_),
    .Y(_1234_));
 sky130_fd_sc_hd__xnor2_1 _2770_ (.A(_0841_),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__a21o_1 _2771_ (.A1(_1227_),
    .A2(_1232_),
    .B1(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__nand3_1 _2772_ (.A(_1227_),
    .B(_1235_),
    .C(_1232_),
    .Y(_1237_));
 sky130_fd_sc_hd__and3_1 _2773_ (.A(_1117_),
    .B(_1236_),
    .C(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2774_ (.A(_1238_),
    .X(_0168_));
 sky130_fd_sc_hd__or3b_1 _2775_ (.A(_1233_),
    .B(_0871_),
    .C_N(_1223_),
    .X(_1239_));
 sky130_fd_sc_hd__inv_2 _2776_ (.A(_0871_),
    .Y(_1240_));
 sky130_fd_sc_hd__a21o_1 _2777_ (.A1(_0854_),
    .A2(_1223_),
    .B1(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__a21oi_1 _2778_ (.A1(_1239_),
    .A2(_1241_),
    .B1(_0858_),
    .Y(_1242_));
 sky130_fd_sc_hd__and3_1 _2779_ (.A(_0858_),
    .B(_1239_),
    .C(_1241_),
    .X(_1243_));
 sky130_fd_sc_hd__nor2_1 _2780_ (.A(_1242_),
    .B(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__or2b_1 _2781_ (.A(_1234_),
    .B_N(_0841_),
    .X(_1245_));
 sky130_fd_sc_hd__nand2_1 _2782_ (.A(_1245_),
    .B(_1237_),
    .Y(_1246_));
 sky130_fd_sc_hd__nand2_1 _2783_ (.A(_1244_),
    .B(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__o211a_1 _2784_ (.A1(_1244_),
    .A2(_1246_),
    .B1(_1247_),
    .C1(_1118_),
    .X(_0169_));
 sky130_fd_sc_hd__and3b_1 _2785_ (.A_N(_1228_),
    .B(_1235_),
    .C(_1244_),
    .X(_1248_));
 sky130_fd_sc_hd__nor2_1 _2786_ (.A(_1245_),
    .B(_1243_),
    .Y(_1249_));
 sky130_fd_sc_hd__a41o_1 _2787_ (.A1(_1227_),
    .A2(_1235_),
    .A3(_1231_),
    .A4(_1244_),
    .B1(_1242_),
    .X(_1250_));
 sky130_fd_sc_hd__a211o_2 _2788_ (.A1(_1220_),
    .A2(_1248_),
    .B1(_1249_),
    .C1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__or4b_1 _2789_ (.A(_0767_),
    .B(_1233_),
    .C(_0871_),
    .D_N(_1223_),
    .X(_1252_));
 sky130_fd_sc_hd__nand2_1 _2790_ (.A(_0767_),
    .B(_1239_),
    .Y(_1253_));
 sky130_fd_sc_hd__a21oi_1 _2791_ (.A1(_1252_),
    .A2(_1253_),
    .B1(_0771_),
    .Y(_1254_));
 sky130_fd_sc_hd__and3_1 _2792_ (.A(_0771_),
    .B(_1252_),
    .C(_1253_),
    .X(_1255_));
 sky130_fd_sc_hd__nor2_1 _2793_ (.A(_1254_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__a21oi_1 _2794_ (.A1(_1251_),
    .A2(_1256_),
    .B1(_1125_),
    .Y(_1257_));
 sky130_fd_sc_hd__o21a_1 _2795_ (.A1(_1251_),
    .A2(_1256_),
    .B1(_1257_),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_1 _2796_ (.A(_0766_),
    .B(_0785_),
    .Y(_1258_));
 sky130_fd_sc_hd__and4_1 _2797_ (.A(_0854_),
    .B(_1240_),
    .C(_1223_),
    .D(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a21o_1 _2798_ (.A1(_0785_),
    .A2(_1252_),
    .B1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__nand2_1 _2799_ (.A(_0789_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__or2_2 _2800_ (.A(_0789_),
    .B(_1260_),
    .X(_1262_));
 sky130_fd_sc_hd__nand2_1 _2801_ (.A(_1261_),
    .B(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__a21oi_1 _2802_ (.A1(_1251_),
    .A2(_1256_),
    .B1(_1254_),
    .Y(_1264_));
 sky130_fd_sc_hd__a21oi_1 _2803_ (.A1(_1263_),
    .A2(_1264_),
    .B1(_1115_),
    .Y(_1265_));
 sky130_fd_sc_hd__o21a_1 _2804_ (.A1(_1263_),
    .A2(_1264_),
    .B1(_1265_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_1 _2805_ (.A(_1261_),
    .B(_1264_),
    .Y(_1266_));
 sky130_fd_sc_hd__inv_2 _2806_ (.A(_0809_),
    .Y(_1267_));
 sky130_fd_sc_hd__xnor2_1 _2807_ (.A(_1267_),
    .B(_1259_),
    .Y(_1268_));
 sky130_fd_sc_hd__xnor2_1 _2808_ (.A(_0796_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__a21oi_1 _2809_ (.A1(_1262_),
    .A2(_1266_),
    .B1(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__a31o_1 _2810_ (.A1(_1262_),
    .A2(_1269_),
    .A3(_1266_),
    .B1(_1115_),
    .X(_1271_));
 sky130_fd_sc_hd__nor2_1 _2811_ (.A(_1270_),
    .B(_1271_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand4_1 _2812_ (.A(_0854_),
    .B(_1240_),
    .C(_1223_),
    .D(_1258_),
    .Y(_1272_));
 sky130_fd_sc_hd__or3_1 _2813_ (.A(_0750_),
    .B(_1267_),
    .C(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__a21o_1 _2814_ (.A1(_0809_),
    .A2(_1259_),
    .B1(_0751_),
    .X(_1274_));
 sky130_fd_sc_hd__and3_1 _2815_ (.A(_0736_),
    .B(_1273_),
    .C(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__a21oi_1 _2816_ (.A1(_1273_),
    .A2(_1274_),
    .B1(_0736_),
    .Y(_1276_));
 sky130_fd_sc_hd__nor2_1 _2817_ (.A(_1275_),
    .B(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__and2b_1 _2818_ (.A_N(_1268_),
    .B(_0796_),
    .X(_1278_));
 sky130_fd_sc_hd__a31o_1 _2819_ (.A1(_1262_),
    .A2(_1269_),
    .A3(_1266_),
    .B1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__nand2_1 _2820_ (.A(_1277_),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__o211a_1 _2821_ (.A1(_1277_),
    .A2(_1279_),
    .B1(_1280_),
    .C1(_1118_),
    .X(_0173_));
 sky130_fd_sc_hd__or4_1 _2822_ (.A(_0731_),
    .B(_0750_),
    .C(_1267_),
    .D(_1272_),
    .X(_1281_));
 sky130_fd_sc_hd__inv_2 _2823_ (.A(_0750_),
    .Y(_1282_));
 sky130_fd_sc_hd__inv_2 _2824_ (.A(_0731_),
    .Y(_1283_));
 sky130_fd_sc_hd__a31o_1 _2825_ (.A1(_1282_),
    .A2(_0809_),
    .A3(_1259_),
    .B1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a21o_1 _2826_ (.A1(_1281_),
    .A2(_1284_),
    .B1(_0717_),
    .X(_1285_));
 sky130_fd_sc_hd__nand3_1 _2827_ (.A(_0717_),
    .B(_1281_),
    .C(_1284_),
    .Y(_1286_));
 sky130_fd_sc_hd__and2_1 _2828_ (.A(_1285_),
    .B(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__and2_1 _2829_ (.A(_0789_),
    .B(_1260_),
    .X(_1288_));
 sky130_fd_sc_hd__or3b_1 _2830_ (.A(_1275_),
    .B(_1276_),
    .C_N(_1269_),
    .X(_1289_));
 sky130_fd_sc_hd__and4bb_1 _2831_ (.A_N(_1288_),
    .B_N(_1289_),
    .C(_1262_),
    .D(_1256_),
    .X(_1290_));
 sky130_fd_sc_hd__o21ai_1 _2832_ (.A1(_1254_),
    .A2(_1288_),
    .B1(_1262_),
    .Y(_1291_));
 sky130_fd_sc_hd__nor2_1 _2833_ (.A(_1278_),
    .B(_1276_),
    .Y(_1292_));
 sky130_fd_sc_hd__o22ai_2 _2834_ (.A1(_1291_),
    .A2(_1289_),
    .B1(_1292_),
    .B2(_1275_),
    .Y(_1293_));
 sky130_fd_sc_hd__a21o_1 _2835_ (.A1(_1251_),
    .A2(_1290_),
    .B1(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__xnor2_1 _2836_ (.A(_1287_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__nor2_1 _2837_ (.A(_1125_),
    .B(_1295_),
    .Y(_0175_));
 sky130_fd_sc_hd__nor2_1 _2838_ (.A(_0712_),
    .B(_0731_),
    .Y(_1296_));
 sky130_fd_sc_hd__and4_1 _2839_ (.A(_1282_),
    .B(_0809_),
    .C(_1259_),
    .D(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_2 _2840_ (.A(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__o41a_1 _2841_ (.A1(_0731_),
    .A2(_0750_),
    .A3(_1267_),
    .A4(_1272_),
    .B1(_0712_),
    .X(_1299_));
 sky130_fd_sc_hd__o21ai_1 _2842_ (.A1(_1298_),
    .A2(_1299_),
    .B1(_0698_),
    .Y(_1300_));
 sky130_fd_sc_hd__or3_1 _2843_ (.A(_0698_),
    .B(_1298_),
    .C(_1299_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _2844_ (.A(_1300_),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__a21boi_1 _2845_ (.A1(_1287_),
    .A2(_1294_),
    .B1_N(_1285_),
    .Y(_1303_));
 sky130_fd_sc_hd__a21oi_1 _2846_ (.A1(_1302_),
    .A2(_1303_),
    .B1(_1115_),
    .Y(_1304_));
 sky130_fd_sc_hd__o21a_1 _2847_ (.A1(_1302_),
    .A2(_1303_),
    .B1(_1304_),
    .X(_0176_));
 sky130_fd_sc_hd__xnor2_1 _2848_ (.A(_0693_),
    .B(_1298_),
    .Y(_1305_));
 sky130_fd_sc_hd__xnor2_1 _2849_ (.A(_0679_),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__a21boi_1 _2850_ (.A1(_1285_),
    .A2(_1300_),
    .B1_N(_1301_),
    .Y(_1307_));
 sky130_fd_sc_hd__a31o_1 _2851_ (.A1(_1287_),
    .A2(_1294_),
    .A3(_1301_),
    .B1(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__xor2_1 _2852_ (.A(_1306_),
    .B(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__nor2_1 _2853_ (.A(_1125_),
    .B(_1309_),
    .Y(_0177_));
 sky130_fd_sc_hd__or3b_1 _2854_ (.A(_0693_),
    .B(_0830_),
    .C_N(_1298_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_2 _2855_ (.A(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__inv_2 _2856_ (.A(_0693_),
    .Y(_1312_));
 sky130_fd_sc_hd__inv_2 _2857_ (.A(_0830_),
    .Y(_1313_));
 sky130_fd_sc_hd__a21o_1 _2858_ (.A1(_1312_),
    .A2(_1298_),
    .B1(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__a21oi_1 _2859_ (.A1(_1311_),
    .A2(_1314_),
    .B1(_0817_),
    .Y(_1315_));
 sky130_fd_sc_hd__nand3_1 _2860_ (.A(_0817_),
    .B(_1311_),
    .C(_1314_),
    .Y(_1316_));
 sky130_fd_sc_hd__and2b_1 _2861_ (.A_N(_1315_),
    .B(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nand2_1 _2862_ (.A(_0679_),
    .B(_1305_),
    .Y(_1318_));
 sky130_fd_sc_hd__nor2_1 _2863_ (.A(_0679_),
    .B(_1305_),
    .Y(_1319_));
 sky130_fd_sc_hd__a21o_1 _2864_ (.A1(_1318_),
    .A2(_1308_),
    .B1(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_1 _2865_ (.A(_1317_),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__o211a_1 _2866_ (.A1(_1317_),
    .A2(_1320_),
    .B1(_1321_),
    .C1(_1118_),
    .X(_0178_));
 sky130_fd_sc_hd__and4_1 _2867_ (.A(_1285_),
    .B(_1286_),
    .C(_1300_),
    .D(_1301_),
    .X(_1322_));
 sky130_fd_sc_hd__and4bb_1 _2868_ (.A_N(_1306_),
    .B_N(_1315_),
    .C(_1316_),
    .D(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__nand3_1 _2869_ (.A(_1251_),
    .B(_1290_),
    .C(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__and4bb_1 _2870_ (.A_N(_1315_),
    .B_N(_1306_),
    .C(_1307_),
    .D(_1316_),
    .X(_1325_));
 sky130_fd_sc_hd__o21a_1 _2871_ (.A1(_1319_),
    .A2(_1315_),
    .B1(_1316_),
    .X(_1326_));
 sky130_fd_sc_hd__a211oi_2 _2872_ (.A1(_1293_),
    .A2(_1323_),
    .B1(_1325_),
    .C1(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__nand2_1 _2873_ (.A(_1324_),
    .B(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_0650_),
    .A1(_0651_),
    .S(_1311_),
    .X(_1329_));
 sky130_fd_sc_hd__xnor2_2 _2875_ (.A(_0637_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__o21ai_1 _2876_ (.A1(_1328_),
    .A2(_1330_),
    .B1(_1117_),
    .Y(_1331_));
 sky130_fd_sc_hd__a21oi_1 _2877_ (.A1(_1328_),
    .A2(_1330_),
    .B1(_1331_),
    .Y(_0179_));
 sky130_fd_sc_hd__nor2_1 _2878_ (.A(_0552_),
    .B(_0650_),
    .Y(_1332_));
 sky130_fd_sc_hd__inv_2 _2879_ (.A(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__inv_2 _2880_ (.A(_0650_),
    .Y(_1334_));
 sky130_fd_sc_hd__a41oi_1 _2881_ (.A1(_1334_),
    .A2(_1312_),
    .A3(_1313_),
    .A4(_1298_),
    .B1(_0553_),
    .Y(_1335_));
 sky130_fd_sc_hd__o21ba_1 _2882_ (.A1(_1311_),
    .A2(_1333_),
    .B1_N(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__xnor2_1 _2883_ (.A(_0535_),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__and2b_1 _2884_ (.A_N(_1329_),
    .B(_0637_),
    .X(_1338_));
 sky130_fd_sc_hd__a21oi_1 _2885_ (.A1(_1328_),
    .A2(_1330_),
    .B1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__xnor2_1 _2886_ (.A(_1337_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__and2_1 _2887_ (.A(_1117_),
    .B(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _2888_ (.A(_1341_),
    .X(_0180_));
 sky130_fd_sc_hd__or3_1 _2889_ (.A(_0570_),
    .B(_1311_),
    .C(_1333_),
    .X(_1342_));
 sky130_fd_sc_hd__o21ai_1 _2890_ (.A1(_1311_),
    .A2(_1333_),
    .B1(_0570_),
    .Y(_1343_));
 sky130_fd_sc_hd__a21oi_1 _2891_ (.A1(_1342_),
    .A2(_1343_),
    .B1(_0557_),
    .Y(_1344_));
 sky130_fd_sc_hd__and3_1 _2892_ (.A(_0557_),
    .B(_1342_),
    .C(_1343_),
    .X(_1345_));
 sky130_fd_sc_hd__nor2_1 _2893_ (.A(_1344_),
    .B(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__nand2_1 _2894_ (.A(_0511_),
    .B(_0534_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _2895_ (.A(_1347_),
    .B(_1336_),
    .Y(_1348_));
 sky130_fd_sc_hd__nor2_1 _2896_ (.A(_1347_),
    .B(_1336_),
    .Y(_1349_));
 sky130_fd_sc_hd__o21a_1 _2897_ (.A1(_1338_),
    .A2(_1349_),
    .B1(_1348_),
    .X(_1350_));
 sky130_fd_sc_hd__a31oi_2 _2898_ (.A1(_1328_),
    .A2(_1330_),
    .A3(_1348_),
    .B1(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__xor2_1 _2899_ (.A(_1346_),
    .B(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__nor2_1 _2900_ (.A(_1125_),
    .B(_1352_),
    .Y(_0181_));
 sky130_fd_sc_hd__or4_2 _2901_ (.A(_0570_),
    .B(_0589_),
    .C(_1311_),
    .D(_1333_),
    .X(_1353_));
 sky130_fd_sc_hd__o31ai_1 _2902_ (.A1(_0570_),
    .A2(_1311_),
    .A3(_1333_),
    .B1(_0591_),
    .Y(_1354_));
 sky130_fd_sc_hd__a21oi_1 _2903_ (.A1(_1353_),
    .A2(_1354_),
    .B1(_0574_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand3_1 _2904_ (.A(_0574_),
    .B(_1353_),
    .C(_1354_),
    .Y(_1356_));
 sky130_fd_sc_hd__and2b_1 _2905_ (.A_N(_1355_),
    .B(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__o21bai_1 _2906_ (.A1(_1345_),
    .A2(_1351_),
    .B1_N(_1344_),
    .Y(_1358_));
 sky130_fd_sc_hd__nand2_1 _2907_ (.A(_1357_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__o211a_1 _2908_ (.A1(_1357_),
    .A2(_1358_),
    .B1(_1359_),
    .C1(_1118_),
    .X(_0182_));
 sky130_fd_sc_hd__or4b_1 _2909_ (.A(_1344_),
    .B(_1345_),
    .C(_1355_),
    .D_N(_1356_),
    .X(_1360_));
 sky130_fd_sc_hd__nand2_1 _2910_ (.A(_1330_),
    .B(_1337_),
    .Y(_1361_));
 sky130_fd_sc_hd__a211o_1 _2911_ (.A1(_1324_),
    .A2(_1327_),
    .B1(_1360_),
    .C1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__o21a_1 _2912_ (.A1(_1344_),
    .A2(_1355_),
    .B1(_1356_),
    .X(_1363_));
 sky130_fd_sc_hd__a31oi_2 _2913_ (.A1(_1346_),
    .A2(_1350_),
    .A3(_1357_),
    .B1(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__xor2_1 _2914_ (.A(_0631_),
    .B(_1353_),
    .X(_1365_));
 sky130_fd_sc_hd__or2_1 _2915_ (.A(_0618_),
    .B(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__nand2_1 _2916_ (.A(_0618_),
    .B(_1365_),
    .Y(_1367_));
 sky130_fd_sc_hd__nand2_1 _2917_ (.A(_1366_),
    .B(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__a21oi_2 _2918_ (.A1(_1362_),
    .A2(_1364_),
    .B1(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__a31o_1 _2919_ (.A1(_1362_),
    .A2(_1364_),
    .A3(_1368_),
    .B1(_1115_),
    .X(_1370_));
 sky130_fd_sc_hd__nor2_1 _2920_ (.A(_1369_),
    .B(_1370_),
    .Y(_0183_));
 sky130_fd_sc_hd__nor2_1 _2921_ (.A(_0618_),
    .B(_1365_),
    .Y(_1371_));
 sky130_fd_sc_hd__nor2_1 _2922_ (.A(_0631_),
    .B(_1353_),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_1 _2923_ (.A(_0613_),
    .B(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__or2_1 _2924_ (.A(_0614_),
    .B(_1372_),
    .X(_1374_));
 sky130_fd_sc_hd__a21o_1 _2925_ (.A1(_1373_),
    .A2(_1374_),
    .B1(_0599_),
    .X(_1375_));
 sky130_fd_sc_hd__nand3_1 _2926_ (.A(_0599_),
    .B(_1373_),
    .C(_1374_),
    .Y(_1376_));
 sky130_fd_sc_hd__o211ai_1 _2927_ (.A1(_1371_),
    .A2(_1369_),
    .B1(_1375_),
    .C1(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__a211o_1 _2928_ (.A1(_1375_),
    .A2(_1376_),
    .B1(_1371_),
    .C1(_1369_),
    .X(_1378_));
 sky130_fd_sc_hd__and3_1 _2929_ (.A(_1117_),
    .B(_1377_),
    .C(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(_1379_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_1 _2931_ (.A(_1366_),
    .B(_1375_),
    .Y(_1380_));
 sky130_fd_sc_hd__inv_2 _2932_ (.A(_0671_),
    .Y(_1381_));
 sky130_fd_sc_hd__xnor2_1 _2933_ (.A(_1381_),
    .B(_1373_),
    .Y(_1382_));
 sky130_fd_sc_hd__xor2_1 _2934_ (.A(_0658_),
    .B(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__o211a_1 _2935_ (.A1(_1369_),
    .A2(_1380_),
    .B1(_1383_),
    .C1(_1376_),
    .X(_1384_));
 sky130_fd_sc_hd__o21a_1 _2936_ (.A1(_1369_),
    .A2(_1380_),
    .B1(_1376_),
    .X(_1385_));
 sky130_fd_sc_hd__o21ai_1 _2937_ (.A1(_1383_),
    .A2(_1385_),
    .B1(_1118_),
    .Y(_1386_));
 sky130_fd_sc_hd__nor2_1 _2938_ (.A(_1384_),
    .B(_1386_),
    .Y(_0186_));
 sky130_fd_sc_hd__and2_1 _2939_ (.A(_0658_),
    .B(_1382_),
    .X(_1387_));
 sky130_fd_sc_hd__nor2_1 _2940_ (.A(_1381_),
    .B(_1373_),
    .Y(_1388_));
 sky130_fd_sc_hd__xnor2_1 _2941_ (.A(_0672_),
    .B(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__or3_1 _2942_ (.A(_1387_),
    .B(_1384_),
    .C(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__o21ai_1 _2943_ (.A1(_1387_),
    .A2(_1384_),
    .B1(_1389_),
    .Y(_1391_));
 sky130_fd_sc_hd__and3_1 _2944_ (.A(_1117_),
    .B(_1390_),
    .C(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _2945_ (.A(_1392_),
    .X(_0187_));
 sky130_fd_sc_hd__inv_2 _2946_ (.A(_0209_),
    .Y(_1393_));
 sky130_fd_sc_hd__or2_1 _2947_ (.A(_0236_),
    .B(_0209_),
    .X(_1394_));
 sky130_fd_sc_hd__o211a_1 _2948_ (.A1(\cpu.INSTRUCTION_EXECUTE_3[7] ),
    .A2(_1393_),
    .B1(_0511_),
    .C1(_1394_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(_0235_),
    .A1(\cpu.INSTRUCTION_EXECUTE_3[8] ),
    .S(_0209_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1395_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_0237_),
    .A1(\cpu.INSTRUCTION_EXECUTE_3[9] ),
    .S(_0209_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _2952_ (.A(_1396_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(_1113_),
    .A1(\cpu.INSTRUCTION_EXECUTE_3[10] ),
    .S(_0209_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_1397_),
    .X(_0205_));
 sky130_fd_sc_hd__o21a_1 _2955_ (.A1(\cpu.INSTRUCTION_EXECUTE_3[7] ),
    .A2(_1393_),
    .B1(_1113_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_1113_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _2957_ (.A(_1398_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1113_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _2959_ (.A(_1399_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _2960_ (.A(_1113_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _2961_ (.A(_1400_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _2962_ (.A(_1113_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_1401_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _2964_ (.A(_1113_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _2965_ (.A(_1402_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _2966_ (.A(_1113_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _2967_ (.A(_1403_),
    .X(_0201_));
 sky130_fd_sc_hd__inv_2 _2968_ (.A(_1000_),
    .Y(\cpu.R2_DATA[0] ));
 sky130_fd_sc_hd__inv_2 _2969_ (.A(_0931_),
    .Y(\cpu.R2_DATA[7] ));
 sky130_fd_sc_hd__buf_4 _2970_ (.A(_0415_),
    .X(_1404_));
 sky130_fd_sc_hd__or2_1 _2971_ (.A(\cpu.INSTRUCTION_DECODE_2[0] ),
    .B(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1405_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(\cpu.INSTRUCTION_DECODE_2[4] ),
    .A1(_0000_),
    .S(_1404_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _2974_ (.A(_1406_),
    .X(_0030_));
 sky130_fd_sc_hd__nor2_4 _2975_ (.A(_0215_),
    .B(_0411_),
    .Y(_1407_));
 sky130_fd_sc_hd__a22o_1 _2976_ (.A1(\cpu.INSTRUCTION_DECODE_2[5] ),
    .A2(_0412_),
    .B1(_0447_),
    .B2(_1407_),
    .X(_0031_));
 sky130_fd_sc_hd__or3b_1 _2977_ (.A(\cpu.PC[4] ),
    .B(\cpu.PC[5] ),
    .C_N(_0216_),
    .X(_1408_));
 sky130_fd_sc_hd__nand2_1 _2978_ (.A(_0446_),
    .B(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__a22o_1 _2979_ (.A1(\cpu.INSTRUCTION_DECODE_2[7] ),
    .A2(_0412_),
    .B1(_1407_),
    .B2(_1409_),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _2980_ (.A(_0216_),
    .B(_0217_),
    .X(_1410_));
 sky130_fd_sc_hd__inv_2 _2981_ (.A(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__o21ba_1 _2982_ (.A1(\cpu.PC[3] ),
    .A2(\cpu.PC[4] ),
    .B1_N(\cpu.PC[5] ),
    .X(_1412_));
 sky130_fd_sc_hd__a21boi_1 _2983_ (.A1(\cpu.PC[4] ),
    .A2(_1411_),
    .B1_N(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__nor2_1 _2984_ (.A(_0206_),
    .B(_0213_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _2985_ (.A(_1414_),
    .B(_0415_),
    .Y(_1415_));
 sky130_fd_sc_hd__buf_4 _2986_ (.A(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__nor2_1 _2987_ (.A(_0446_),
    .B(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__a221o_1 _2988_ (.A1(\cpu.INSTRUCTION_DECODE_2[9] ),
    .A2(_0412_),
    .B1(_1407_),
    .B2(_1413_),
    .C1(_1417_),
    .X(_0033_));
 sky130_fd_sc_hd__a31o_1 _2989_ (.A1(\cpu.PC[4] ),
    .A2(_0217_),
    .A3(_1414_),
    .B1(_0004_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(\cpu.INSTRUCTION_DECODE_2[16] ),
    .A1(_0040_),
    .S(_1404_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _2991_ (.A(_1418_),
    .X(_0034_));
 sky130_fd_sc_hd__or3b_1 _2992_ (.A(\cpu.PC[2] ),
    .B(\cpu.PC[5] ),
    .C_N(\cpu.PC[3] ),
    .X(_1419_));
 sky130_fd_sc_hd__a21oi_1 _2993_ (.A1(_1408_),
    .A2(_1419_),
    .B1(_0215_),
    .Y(_0145_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(\cpu.INSTRUCTION_DECODE_2[20] ),
    .A1(_0145_),
    .S(_1404_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _2995_ (.A(_1420_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(\cpu.INSTRUCTION_DECODE_2[21] ),
    .A1(_0002_),
    .S(_1404_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _2997_ (.A(_1421_),
    .X(_0036_));
 sky130_fd_sc_hd__a31o_1 _2998_ (.A1(_1411_),
    .A2(_1414_),
    .A3(_1412_),
    .B1(_0004_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(\cpu.INSTRUCTION_DECODE_2[22] ),
    .A1(_0147_),
    .S(_1404_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _3000_ (.A(_1422_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(\cpu.INSTRUCTION_DECODE_2[11] ),
    .A1(_0004_),
    .S(_1404_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _3002_ (.A(_1423_),
    .X(_0038_));
 sky130_fd_sc_hd__o2bb2ai_1 _3003_ (.A1_N(\cpu.INSTRUCTION_DECODE_2[13] ),
    .A2_N(_0412_),
    .B1(_1416_),
    .B2(_0218_),
    .Y(_0039_));
 sky130_fd_sc_hd__a21oi_1 _3004_ (.A1(\cpu.PC[4] ),
    .A2(_0216_),
    .B1(_0217_),
    .Y(_1424_));
 sky130_fd_sc_hd__inv_2 _3005_ (.A(\cpu.INSTRUCTION_DECODE_2[8] ),
    .Y(_1425_));
 sky130_fd_sc_hd__o32a_1 _3006_ (.A1(\cpu.PC[5] ),
    .A2(_1416_),
    .A3(_1424_),
    .B1(_1425_),
    .B2(_0420_),
    .X(_1426_));
 sky130_fd_sc_hd__clkinv_2 _3007_ (.A(_1426_),
    .Y(_0041_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(\cpu.PC_EXECUTE_3[0] ),
    .A1(\cpu.PC_DECODE_2[0] ),
    .S(_1404_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _3009_ (.A(_1427_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(\cpu.PC_EXECUTE_3[1] ),
    .A1(\cpu.PC_DECODE_2[1] ),
    .S(_1404_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_1428_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(\cpu.PC_EXECUTE_3[2] ),
    .A1(\cpu.PC_DECODE_2[2] ),
    .S(_1404_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _3013_ (.A(_1429_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(\cpu.PC_EXECUTE_3[3] ),
    .A1(\cpu.PC_DECODE_2[3] ),
    .S(_0416_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _3015_ (.A(_1430_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(\cpu.PC_EXECUTE_3[4] ),
    .A1(\cpu.PC_DECODE_2[4] ),
    .S(_0416_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _3017_ (.A(_1431_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(\cpu.PC_EXECUTE_3[5] ),
    .A1(\cpu.PC_DECODE_2[5] ),
    .S(_0416_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1432_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(\cpu.PC_EXECUTE_3[6] ),
    .A1(\cpu.PC_DECODE_2[6] ),
    .S(_0416_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_1433_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(\cpu.PC_EXECUTE_3[7] ),
    .A1(\cpu.PC_DECODE_2[7] ),
    .S(_0416_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3023_ (.A(_1434_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(\cpu.PC_EXECUTE_3[8] ),
    .A1(\cpu.PC_DECODE_2[8] ),
    .S(_0416_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3025_ (.A(_1435_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(\cpu.PC_EXECUTE_3[9] ),
    .A1(\cpu.PC_DECODE_2[9] ),
    .S(_0416_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _3027_ (.A(_1436_),
    .X(_0051_));
 sky130_fd_sc_hd__or4_1 _3028_ (.A(\cpu.ALU_OUT[23] ),
    .B(\cpu.ALU_OUT[22] ),
    .C(\cpu.ALU_OUT[24] ),
    .D(\cpu.ALU_OUT[29] ),
    .X(_1437_));
 sky130_fd_sc_hd__or4_1 _3029_ (.A(\cpu.ALU_OUT[20] ),
    .B(\cpu.ALU_OUT[25] ),
    .C(\cpu.ALU_OUT[27] ),
    .D(\cpu.ALU_OUT[26] ),
    .X(_1438_));
 sky130_fd_sc_hd__or4_2 _3030_ (.A(\cpu.ALU_OUT[28] ),
    .B(\cpu.ALU_OUT[31] ),
    .C(\cpu.ALU_OUT[30] ),
    .D(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__or4_1 _3031_ (.A(\cpu.ALU_OUT[0] ),
    .B(\cpu.ALU_OUT[3] ),
    .C(\cpu.ALU_OUT[2] ),
    .D(\cpu.ALU_OUT[5] ),
    .X(_1440_));
 sky130_fd_sc_hd__or3b_2 _3032_ (.A(\cpu.ALU_OUT[1] ),
    .B(_1440_),
    .C_N(\cpu.TYPE_PIPELINE[1][2] ),
    .X(_1441_));
 sky130_fd_sc_hd__or4_1 _3033_ (.A(\cpu.ALU_OUT[12] ),
    .B(\cpu.ALU_OUT[15] ),
    .C(\cpu.ALU_OUT[14] ),
    .D(\cpu.ALU_OUT[17] ),
    .X(_1442_));
 sky130_fd_sc_hd__or4_1 _3034_ (.A(\cpu.ALU_OUT[8] ),
    .B(\cpu.ALU_OUT[11] ),
    .C(\cpu.ALU_OUT[10] ),
    .D(\cpu.ALU_OUT[13] ),
    .X(_1443_));
 sky130_fd_sc_hd__or4_2 _3035_ (.A(\cpu.ALU_OUT[4] ),
    .B(\cpu.ALU_OUT[7] ),
    .C(\cpu.ALU_OUT[6] ),
    .D(\cpu.ALU_OUT[9] ),
    .X(_1444_));
 sky130_fd_sc_hd__or4_1 _3036_ (.A(\cpu.ALU_OUT[16] ),
    .B(\cpu.ALU_OUT[19] ),
    .C(\cpu.ALU_OUT[18] ),
    .D(\cpu.ALU_OUT[21] ),
    .X(_1445_));
 sky130_fd_sc_hd__or3_1 _3037_ (.A(_1443_),
    .B(_1444_),
    .C(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__or3_2 _3038_ (.A(_1441_),
    .B(_1442_),
    .C(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__nor3_4 _3039_ (.A(_1437_),
    .B(_1439_),
    .C(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__buf_6 _3040_ (.A(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(net1),
    .A1(\cpu.R2_DATA[0] ),
    .S(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3042_ (.A(_1450_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(net12),
    .A1(\cpu.R2_DATA[1] ),
    .S(_1449_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _3044_ (.A(_1451_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(net23),
    .A1(\cpu.R2_DATA[2] ),
    .S(_1449_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1452_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(net26),
    .A1(\cpu.R2_DATA[3] ),
    .S(_1449_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _3048_ (.A(_1453_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(net27),
    .A1(\cpu.R2_DATA[4] ),
    .S(_1449_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _3050_ (.A(_1454_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(net28),
    .A1(\cpu.R2_DATA[5] ),
    .S(_1449_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _3052_ (.A(_1455_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(net29),
    .A1(\cpu.R2_DATA[6] ),
    .S(_1449_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _3054_ (.A(_1456_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(net30),
    .A1(\cpu.R2_DATA[7] ),
    .S(_1449_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3056_ (.A(_1457_),
    .X(_0059_));
 sky130_fd_sc_hd__inv_2 _3057_ (.A(_0950_),
    .Y(_1458_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(net31),
    .A1(_1458_),
    .S(_1449_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _3059_ (.A(_1459_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _3060_ (.A(_1047_),
    .Y(_1460_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(net32),
    .A1(_1460_),
    .S(_1449_),
    .X(_1461_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1461_),
    .X(_0061_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(_1066_),
    .Y(_1462_));
 sky130_fd_sc_hd__buf_6 _3064_ (.A(_1448_),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(net2),
    .A1(_1462_),
    .S(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1464_),
    .X(_0062_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(_1085_),
    .Y(_1465_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(net3),
    .A1(_1465_),
    .S(_1463_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _3069_ (.A(_1466_),
    .X(_0063_));
 sky130_fd_sc_hd__inv_2 _3070_ (.A(_0910_),
    .Y(_1467_));
 sky130_fd_sc_hd__mux2_1 _3071_ (.A0(net4),
    .A1(_1467_),
    .S(_1463_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _3072_ (.A(_1468_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(net5),
    .A1(_0891_),
    .S(_1463_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3074_ (.A(_1469_),
    .X(_0065_));
 sky130_fd_sc_hd__inv_2 _3075_ (.A(_0853_),
    .Y(_1470_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(net6),
    .A1(_1470_),
    .S(_1463_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3077_ (.A(_1471_),
    .X(_0066_));
 sky130_fd_sc_hd__inv_2 _3078_ (.A(_0870_),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(net7),
    .A1(_1472_),
    .S(_1463_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1473_),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _3081_ (.A(_0765_),
    .Y(_1474_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(net8),
    .A1(_1474_),
    .S(_1463_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _3083_ (.A(_1475_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(net9),
    .A1(_0784_),
    .S(_1463_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3085_ (.A(_1476_),
    .X(_0069_));
 sky130_fd_sc_hd__inv_2 _3086_ (.A(_0808_),
    .Y(_1477_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(net10),
    .A1(_1477_),
    .S(_1463_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3088_ (.A(_1478_),
    .X(_0070_));
 sky130_fd_sc_hd__inv_2 _3089_ (.A(_0749_),
    .Y(_1479_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(net11),
    .A1(_1479_),
    .S(_1463_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3091_ (.A(_1480_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_8 _3092_ (.A(_1448_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(net13),
    .A1(_0730_),
    .S(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__clkbuf_1 _3094_ (.A(_1482_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(net14),
    .A1(_0711_),
    .S(_1481_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3096_ (.A(_1483_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(net15),
    .A1(_0692_),
    .S(_1481_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1484_),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _3099_ (.A(_0829_),
    .Y(_1485_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(net16),
    .A1(_1485_),
    .S(_1481_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3101_ (.A(_1486_),
    .X(_0075_));
 sky130_fd_sc_hd__inv_2 _3102_ (.A(_0649_),
    .Y(_1487_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(net17),
    .A1(_1487_),
    .S(_1481_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_1 _3104_ (.A(_1488_),
    .X(_0076_));
 sky130_fd_sc_hd__inv_2 _3105_ (.A(_0549_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(net18),
    .A1(_1489_),
    .S(_1481_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3107_ (.A(_1490_),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _3108_ (.A(_0569_),
    .Y(_1491_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(net19),
    .A1(_1491_),
    .S(_1481_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_1 _3110_ (.A(_1492_),
    .X(_0078_));
 sky130_fd_sc_hd__inv_2 _3111_ (.A(_0588_),
    .Y(_1493_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(net20),
    .A1(_1493_),
    .S(_1481_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_1 _3113_ (.A(_1494_),
    .X(_0079_));
 sky130_fd_sc_hd__inv_2 _3114_ (.A(_0630_),
    .Y(_1495_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(net21),
    .A1(_1495_),
    .S(_1481_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3116_ (.A(_1496_),
    .X(_0080_));
 sky130_fd_sc_hd__inv_2 _3117_ (.A(_0612_),
    .Y(_1497_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(net22),
    .A1(_1497_),
    .S(_1481_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3119_ (.A(_1498_),
    .X(_0081_));
 sky130_fd_sc_hd__inv_2 _3120_ (.A(_0670_),
    .Y(_1499_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(net24),
    .A1(_1499_),
    .S(_1448_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3122_ (.A(_1500_),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _3123_ (.A(_0504_),
    .Y(_1501_));
 sky130_fd_sc_hd__mux2_1 _3124_ (.A0(net25),
    .A1(_1501_),
    .S(_1448_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _3125_ (.A(_1502_),
    .X(_0083_));
 sky130_fd_sc_hd__inv_2 _3126_ (.A(_0975_),
    .Y(_1503_));
 sky130_fd_sc_hd__a211o_1 _3127_ (.A1(_0285_),
    .A2(_0982_),
    .B1(_1000_),
    .C1(_1005_),
    .X(_1504_));
 sky130_fd_sc_hd__a21o_1 _3128_ (.A1(_0328_),
    .A2(_0329_),
    .B1(_1011_),
    .X(_1505_));
 sky130_fd_sc_hd__o211a_1 _3129_ (.A1(_0285_),
    .A2(_0982_),
    .B1(_1504_),
    .C1(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__and3_1 _3130_ (.A(_0328_),
    .B(_0329_),
    .C(_1011_),
    .X(_1507_));
 sky130_fd_sc_hd__and3_1 _3131_ (.A(_0288_),
    .B(_0312_),
    .C(_1019_),
    .X(_1508_));
 sky130_fd_sc_hd__a21o_1 _3132_ (.A1(_0288_),
    .A2(_0312_),
    .B1(_1019_),
    .X(_1509_));
 sky130_fd_sc_hd__nand2_1 _3133_ (.A(\cpu.R2_DATA[4] ),
    .B(_1503_),
    .Y(_1510_));
 sky130_fd_sc_hd__o311ai_1 _3134_ (.A1(_1506_),
    .A2(_1507_),
    .A3(_1508_),
    .B1(_1509_),
    .C1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__o221a_1 _3135_ (.A1(\cpu.R2_DATA[5] ),
    .A2(_0960_),
    .B1(_1503_),
    .B2(\cpu.R2_DATA[4] ),
    .C1(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__a221o_1 _3136_ (.A1(\cpu.R2_DATA[6] ),
    .A2(_0966_),
    .B1(_0960_),
    .B2(\cpu.R2_DATA[5] ),
    .C1(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__o2bb2a_1 _3137_ (.A1_N(_0931_),
    .A2_N(_0917_),
    .B1(_0966_),
    .B2(\cpu.R2_DATA[6] ),
    .X(_1514_));
 sky130_fd_sc_hd__o22ai_1 _3138_ (.A1(_0950_),
    .A2(_0936_),
    .B1(_0931_),
    .B2(_0917_),
    .Y(_1515_));
 sky130_fd_sc_hd__a21oi_1 _3139_ (.A1(_1513_),
    .A2(_1514_),
    .B1(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__a221o_1 _3140_ (.A1(_0950_),
    .A2(_0936_),
    .B1(_1047_),
    .B2(_1033_),
    .C1(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__o22a_1 _3141_ (.A1(_1053_),
    .A2(_1066_),
    .B1(_1047_),
    .B2(_1033_),
    .X(_1518_));
 sky130_fd_sc_hd__a22o_1 _3142_ (.A1(_1053_),
    .A2(_1066_),
    .B1(_1071_),
    .B2(_1085_),
    .X(_1519_));
 sky130_fd_sc_hd__a21oi_1 _3143_ (.A1(_1517_),
    .A2(_1518_),
    .B1(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__a22o_1 _3144_ (.A1(_0840_),
    .A2(_0853_),
    .B1(_0857_),
    .B2(_0870_),
    .X(_1521_));
 sky130_fd_sc_hd__or2_1 _3145_ (.A(_0857_),
    .B(_0870_),
    .X(_1522_));
 sky130_fd_sc_hd__o221a_1 _3146_ (.A1(_0840_),
    .A2(_0853_),
    .B1(_0877_),
    .B2(_0890_),
    .C1(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__or2b_1 _3147_ (.A(_1521_),
    .B_N(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__a22oi_1 _3148_ (.A1(_0877_),
    .A2(_0890_),
    .B1(_0897_),
    .B2(_0910_),
    .Y(_1525_));
 sky130_fd_sc_hd__o221ai_1 _3149_ (.A1(_1071_),
    .A2(_1085_),
    .B1(_0897_),
    .B2(_0910_),
    .C1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__o2bb2a_1 _3150_ (.A1_N(_1521_),
    .A2_N(_1522_),
    .B1(_1524_),
    .B2(_1525_),
    .X(_1527_));
 sky130_fd_sc_hd__o31a_1 _3151_ (.A1(_1520_),
    .A2(_1524_),
    .A3(_1526_),
    .B1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__o21ai_1 _3152_ (.A1(\cpu.ALU_OUT_MEMORY_4[21] ),
    .A2(_0451_),
    .B1(_0710_),
    .Y(_1529_));
 sky130_fd_sc_hd__a22o_1 _3153_ (.A1(_0697_),
    .A2(_1529_),
    .B1(_0716_),
    .B2(_0729_),
    .X(_1530_));
 sky130_fd_sc_hd__o22ai_1 _3154_ (.A1(_0678_),
    .A2(_0691_),
    .B1(_0697_),
    .B2(_1529_),
    .Y(_1531_));
 sky130_fd_sc_hd__or2_1 _3155_ (.A(_0716_),
    .B(_0729_),
    .X(_1532_));
 sky130_fd_sc_hd__or2_1 _3156_ (.A(_0795_),
    .B(_0808_),
    .X(_1533_));
 sky130_fd_sc_hd__or2_1 _3157_ (.A(_0783_),
    .B(_0788_),
    .X(_1534_));
 sky130_fd_sc_hd__or2_1 _3158_ (.A(_0735_),
    .B(_0749_),
    .X(_1535_));
 sky130_fd_sc_hd__and3_1 _3159_ (.A(_1533_),
    .B(_1534_),
    .C(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__o211a_1 _3160_ (.A1(_0765_),
    .A2(_0770_),
    .B1(_1532_),
    .C1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__or3b_1 _3161_ (.A(_1530_),
    .B(_1531_),
    .C_N(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__a22o_1 _3162_ (.A1(_0678_),
    .A2(_0691_),
    .B1(_0816_),
    .B2(_0829_),
    .X(_1539_));
 sky130_fd_sc_hd__a22o_1 _3163_ (.A1(_0735_),
    .A2(_0749_),
    .B1(_0795_),
    .B2(_0808_),
    .X(_1540_));
 sky130_fd_sc_hd__a22o_1 _3164_ (.A1(_0765_),
    .A2(_0770_),
    .B1(_0783_),
    .B2(_0788_),
    .X(_1541_));
 sky130_fd_sc_hd__or2_1 _3165_ (.A(_0816_),
    .B(_0829_),
    .X(_1542_));
 sky130_fd_sc_hd__or4b_1 _3166_ (.A(_1539_),
    .B(_1540_),
    .C(_1541_),
    .D_N(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__a31o_1 _3167_ (.A1(_1541_),
    .A2(_1533_),
    .A3(_1534_),
    .B1(_1540_),
    .X(_1544_));
 sky130_fd_sc_hd__a31o_1 _3168_ (.A1(_1544_),
    .A2(_1532_),
    .A3(_1535_),
    .B1(_1530_),
    .X(_1545_));
 sky130_fd_sc_hd__and2b_1 _3169_ (.A_N(_1531_),
    .B(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__o21ai_1 _3170_ (.A1(_1539_),
    .A2(_1546_),
    .B1(_1542_),
    .Y(_1547_));
 sky130_fd_sc_hd__o31a_1 _3171_ (.A1(_1528_),
    .A2(_1538_),
    .A3(_1543_),
    .B1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__o22a_1 _3172_ (.A1(_0556_),
    .A2(_0569_),
    .B1(_0534_),
    .B2(_0549_),
    .X(_1549_));
 sky130_fd_sc_hd__a22o_1 _3173_ (.A1(_0556_),
    .A2(_0569_),
    .B1(_0573_),
    .B2(_0588_),
    .X(_1550_));
 sky130_fd_sc_hd__a22o_1 _3174_ (.A1(_0534_),
    .A2(_0549_),
    .B1(_0636_),
    .B2(_0649_),
    .X(_1551_));
 sky130_fd_sc_hd__nor2_1 _3175_ (.A(_1550_),
    .B(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__a22o_1 _3176_ (.A1(_0598_),
    .A2(_0612_),
    .B1(_0617_),
    .B2(_0630_),
    .X(_1553_));
 sky130_fd_sc_hd__o22ai_1 _3177_ (.A1(_0573_),
    .A2(_0588_),
    .B1(_0617_),
    .B2(_0630_),
    .Y(_1554_));
 sky130_fd_sc_hd__nor2_1 _3178_ (.A(_1553_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__xor2_2 _3179_ (.A(_0529_),
    .B(_0504_),
    .X(_1556_));
 sky130_fd_sc_hd__o22ai_1 _3180_ (.A1(_0657_),
    .A2(_0670_),
    .B1(_0598_),
    .B2(_0612_),
    .Y(_1557_));
 sky130_fd_sc_hd__and2_1 _3181_ (.A(_0657_),
    .B(_0670_),
    .X(_1558_));
 sky130_fd_sc_hd__nor2_1 _3182_ (.A(_1557_),
    .B(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__o2111a_1 _3183_ (.A1(_0636_),
    .A2(_0649_),
    .B1(_1555_),
    .C1(_1556_),
    .D1(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__and4b_1 _3184_ (.A_N(_1548_),
    .B(_1549_),
    .C(_1552_),
    .D(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__a21oi_1 _3185_ (.A1(_1549_),
    .A2(_1551_),
    .B1(_1550_),
    .Y(_1562_));
 sky130_fd_sc_hd__nor2_1 _3186_ (.A(_1554_),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__o21ba_1 _3187_ (.A1(_1553_),
    .A2(_1563_),
    .B1_N(_1557_),
    .X(_1564_));
 sky130_fd_sc_hd__o22a_1 _3188_ (.A1(_0529_),
    .A2(_0504_),
    .B1(_1558_),
    .B2(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__a211o_2 _3189_ (.A1(_0529_),
    .A2(_0504_),
    .B1(_1561_),
    .C1(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__or2_1 _3190_ (.A(\cpu.INSTRUCTION_EXECUTE_3[13] ),
    .B(_1556_),
    .X(_1567_));
 sky130_fd_sc_hd__a21oi_1 _3191_ (.A1(_1566_),
    .A2(_1567_),
    .B1(_0511_),
    .Y(_1568_));
 sky130_fd_sc_hd__o21ai_4 _3192_ (.A1(_1566_),
    .A2(_1567_),
    .B1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\cpu.ALU_OUT[0] ),
    .A1(\cpu.PC[0] ),
    .S(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_1570_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(\cpu.ALU_OUT[1] ),
    .A1(\cpu.PC[1] ),
    .S(_1569_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3196_ (.A(_1571_),
    .X(_0085_));
 sky130_fd_sc_hd__and3_1 _3197_ (.A(\cpu.PC[2] ),
    .B(\cpu.PC[3] ),
    .C(_1407_),
    .X(_1572_));
 sky130_fd_sc_hd__a22o_1 _3198_ (.A1(\cpu.INSTRUCTION_DECODE_2[10] ),
    .A2(_0412_),
    .B1(_1413_),
    .B2(_1572_),
    .X(_0086_));
 sky130_fd_sc_hd__buf_4 _3199_ (.A(_0422_),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(\cpu.ALU_OUT_MEMORY_4[11] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[11] ),
    .S(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _3201_ (.A(_1574_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(\cpu.ALU_OUT_MEMORY_4[12] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[12] ),
    .S(_1573_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_1575_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(\cpu.ALU_OUT_MEMORY_4[13] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[13] ),
    .S(_1573_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3205_ (.A(_1576_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(\cpu.ALU_OUT_MEMORY_4[14] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[14] ),
    .S(_1573_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _3207_ (.A(_1577_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(\cpu.ALU_OUT_MEMORY_4[15] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[15] ),
    .S(_1573_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _3209_ (.A(_1578_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(\cpu.ALU_OUT_MEMORY_4[16] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[16] ),
    .S(_1573_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3211_ (.A(_1579_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(\cpu.ALU_OUT_MEMORY_4[17] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[17] ),
    .S(_1573_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3213_ (.A(_1580_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(\cpu.ALU_OUT_MEMORY_4[18] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[18] ),
    .S(_1573_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3215_ (.A(_1581_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(\cpu.ALU_OUT_MEMORY_4[19] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[19] ),
    .S(_1573_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3217_ (.A(_1582_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(\cpu.ALU_OUT_MEMORY_4[20] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[20] ),
    .S(_1573_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_1583_),
    .X(_0096_));
 sky130_fd_sc_hd__buf_4 _3220_ (.A(_0422_),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\cpu.ALU_OUT_MEMORY_4[21] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[21] ),
    .S(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3222_ (.A(_1585_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\cpu.ALU_OUT_MEMORY_4[22] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[22] ),
    .S(_1584_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3224_ (.A(_1586_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(\cpu.ALU_OUT_MEMORY_4[23] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[23] ),
    .S(_1584_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1587_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\cpu.ALU_OUT_MEMORY_4[24] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[24] ),
    .S(_1584_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _3228_ (.A(_1588_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(\cpu.ALU_OUT_MEMORY_4[25] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[25] ),
    .S(_1584_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3230_ (.A(_1589_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(\cpu.ALU_OUT_MEMORY_4[26] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[26] ),
    .S(_1584_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_1590_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(\cpu.ALU_OUT_MEMORY_4[27] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[27] ),
    .S(_1584_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3234_ (.A(_1591_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(\cpu.ALU_OUT_MEMORY_4[28] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[28] ),
    .S(_1584_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _3236_ (.A(_1592_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(\cpu.ALU_OUT_MEMORY_4[29] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[29] ),
    .S(_1584_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_1593_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(\cpu.ALU_OUT_MEMORY_4[30] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[30] ),
    .S(_1584_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3240_ (.A(_1594_),
    .X(_0106_));
 sky130_fd_sc_hd__buf_6 _3241_ (.A(_0422_),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(\cpu.ALU_OUT_MEMORY_4[31] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[31] ),
    .S(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3243_ (.A(_1596_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(\cpu.PC_DECODE_2[0] ),
    .A1(\cpu.PC[0] ),
    .S(_1407_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3245_ (.A(_1597_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(\cpu.PC_DECODE_2[1] ),
    .A1(\cpu.PC[1] ),
    .S(_1407_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_1598_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(\cpu.PC[2] ),
    .A1(\cpu.PC_DECODE_2[2] ),
    .S(_1416_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _3249_ (.A(_1599_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(\cpu.PC[3] ),
    .A1(\cpu.PC_DECODE_2[3] ),
    .S(_1416_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3251_ (.A(_1600_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(\cpu.PC[4] ),
    .A1(\cpu.PC_DECODE_2[4] ),
    .S(_1416_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_1601_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(\cpu.PC[5] ),
    .A1(\cpu.PC_DECODE_2[5] ),
    .S(_1416_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1602_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(\cpu.PC[6] ),
    .A1(\cpu.PC_DECODE_2[6] ),
    .S(_1416_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _3257_ (.A(_1603_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(\cpu.PC[7] ),
    .A1(\cpu.PC_DECODE_2[7] ),
    .S(_1416_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_1604_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(\cpu.PC[8] ),
    .A1(\cpu.PC_DECODE_2[8] ),
    .S(_1416_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3261_ (.A(_1605_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\cpu.PC[9] ),
    .A1(\cpu.PC_DECODE_2[9] ),
    .S(_1415_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3263_ (.A(_1606_),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _3264_ (.A(\cpu.INSTRUCTION_DECODE_2[0] ),
    .B(_0412_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_1607_),
    .X(_0118_));
 sky130_fd_sc_hd__nand2_1 _3266_ (.A(_0212_),
    .B(_0420_),
    .Y(_0119_));
 sky130_fd_sc_hd__and2_1 _3267_ (.A(\cpu.INSTRUCTION_DECODE_2[7] ),
    .B(_0420_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3268_ (.A(_1608_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _3269_ (.A(_1425_),
    .B(_0412_),
    .Y(_0122_));
 sky130_fd_sc_hd__and2_1 _3270_ (.A(\cpu.INSTRUCTION_DECODE_2[9] ),
    .B(_0420_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_1 _3271_ (.A(_1609_),
    .X(_0123_));
 sky130_fd_sc_hd__and2_1 _3272_ (.A(\cpu.INSTRUCTION_DECODE_2[10] ),
    .B(_0420_),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1610_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _3274_ (.A(\cpu.INSTRUCTION_DECODE_2[13] ),
    .B(_0420_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3275_ (.A(_1611_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _3276_ (.A(\cpu.INSTRUCTION_DECODE_2[16] ),
    .B(_0420_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _3277_ (.A(_1612_),
    .X(_0126_));
 sky130_fd_sc_hd__and2_1 _3278_ (.A(\cpu.INSTRUCTION_DECODE_2[20] ),
    .B(_0420_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_1 _3279_ (.A(_1613_),
    .X(_0127_));
 sky130_fd_sc_hd__and2_1 _3280_ (.A(\cpu.INSTRUCTION_DECODE_2[21] ),
    .B(_0420_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _3281_ (.A(_1614_),
    .X(_0128_));
 sky130_fd_sc_hd__buf_2 _3282_ (.A(_0416_),
    .X(_1615_));
 sky130_fd_sc_hd__and2_1 _3283_ (.A(\cpu.INSTRUCTION_DECODE_2[22] ),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3284_ (.A(_1616_),
    .X(_0129_));
 sky130_fd_sc_hd__and2_1 _3285_ (.A(\cpu.INSTRUCTION_DECODE_2[11] ),
    .B(_1615_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3286_ (.A(_1617_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _3287_ (.A(\cpu.INSTRUCTION_DECODE_2[16] ),
    .B(_1615_),
    .X(_1618_));
 sky130_fd_sc_hd__clkbuf_1 _3288_ (.A(_1618_),
    .X(_0131_));
 sky130_fd_sc_hd__xnor2_1 _3289_ (.A(\cpu.PC[2] ),
    .B(_1415_),
    .Y(_1619_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\cpu.ALU_OUT[2] ),
    .A1(_1619_),
    .S(_1569_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1620_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\cpu.PC[3] ),
    .A1(_1410_),
    .S(_1407_),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(\cpu.ALU_OUT[3] ),
    .A1(_1621_),
    .S(_1569_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _3294_ (.A(_1622_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _3295_ (.A(\cpu.PC[4] ),
    .B(_1572_),
    .X(_1623_));
 sky130_fd_sc_hd__nor2_1 _3296_ (.A(\cpu.PC[4] ),
    .B(_1572_),
    .Y(_1624_));
 sky130_fd_sc_hd__nor2_1 _3297_ (.A(_1623_),
    .B(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(\cpu.ALU_OUT[4] ),
    .A1(_1625_),
    .S(_1569_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _3299_ (.A(_1626_),
    .X(_0134_));
 sky130_fd_sc_hd__xor2_1 _3300_ (.A(\cpu.PC[5] ),
    .B(_1623_),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(\cpu.ALU_OUT[5] ),
    .A1(_1627_),
    .S(_1569_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _3302_ (.A(_1628_),
    .X(_0135_));
 sky130_fd_sc_hd__and3_1 _3303_ (.A(\cpu.PC[5] ),
    .B(\cpu.PC[6] ),
    .C(_1623_),
    .X(_1629_));
 sky130_fd_sc_hd__a21oi_1 _3304_ (.A1(\cpu.PC[5] ),
    .A2(_1623_),
    .B1(\cpu.PC[6] ),
    .Y(_1630_));
 sky130_fd_sc_hd__nor2_1 _3305_ (.A(_1629_),
    .B(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(\cpu.ALU_OUT[6] ),
    .A1(_1631_),
    .S(_1569_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _3307_ (.A(_1632_),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _3308_ (.A(\cpu.PC[7] ),
    .B(_1629_),
    .X(_1633_));
 sky130_fd_sc_hd__nor2_1 _3309_ (.A(\cpu.PC[7] ),
    .B(_1629_),
    .Y(_1634_));
 sky130_fd_sc_hd__nor2_1 _3310_ (.A(_1633_),
    .B(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(\cpu.ALU_OUT[7] ),
    .A1(_1635_),
    .S(_1569_),
    .X(_1636_));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(_1636_),
    .X(_0137_));
 sky130_fd_sc_hd__nand2_1 _3313_ (.A(\cpu.PC[8] ),
    .B(_1633_),
    .Y(_1637_));
 sky130_fd_sc_hd__or2_1 _3314_ (.A(\cpu.PC[8] ),
    .B(_1633_),
    .X(_1638_));
 sky130_fd_sc_hd__and2_1 _3315_ (.A(_1637_),
    .B(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(\cpu.ALU_OUT[8] ),
    .A1(_1639_),
    .S(_1569_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3317_ (.A(_1640_),
    .X(_0138_));
 sky130_fd_sc_hd__xnor2_1 _3318_ (.A(\cpu.PC[9] ),
    .B(_1637_),
    .Y(_1641_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(\cpu.ALU_OUT[9] ),
    .A1(_1641_),
    .S(_1569_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _3320_ (.A(_1642_),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _3321_ (.A(\cpu.INSTRUCTION_DECODE_2[7] ),
    .B(_1615_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _3322_ (.A(_1643_),
    .X(_0140_));
 sky130_fd_sc_hd__nor2_1 _3323_ (.A(_1425_),
    .B(_0412_),
    .Y(_0141_));
 sky130_fd_sc_hd__and2_1 _3324_ (.A(\cpu.INSTRUCTION_DECODE_2[9] ),
    .B(_1615_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _3325_ (.A(_1644_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_1 _3326_ (.A(\cpu.INSTRUCTION_DECODE_2[10] ),
    .B(_1615_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3327_ (.A(_1645_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _3328_ (.A(\cpu.INSTRUCTION_DECODE_2[11] ),
    .B(_1615_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _3329_ (.A(_1646_),
    .X(_0144_));
 sky130_fd_sc_hd__nor2_1 _3330_ (.A(_0215_),
    .B(_0219_),
    .Y(_0146_));
 sky130_fd_sc_hd__nor2_1 _3331_ (.A(_0215_),
    .B(_0446_),
    .Y(_0148_));
 sky130_fd_sc_hd__and2_1 _3332_ (.A(\cpu.INSTRUCTION_DECODE_2[20] ),
    .B(_1615_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3333_ (.A(_1647_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _3334_ (.A(\cpu.INSTRUCTION_DECODE_2[21] ),
    .B(_1615_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _3335_ (.A(_1648_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_1 _3336_ (.A(\cpu.INSTRUCTION_DECODE_2[22] ),
    .B(_1615_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _3337_ (.A(_1649_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _3338_ (.A0(net216),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[0] ),
    .S(_1595_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _3339_ (.A(_1650_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(net210),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[1] ),
    .S(_1595_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _3341_ (.A(_1651_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(net204),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[2] ),
    .S(_1595_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _3343_ (.A(_1652_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(net199),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[3] ),
    .S(_1595_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _3345_ (.A(_1653_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(net193),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[4] ),
    .S(_1595_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3347_ (.A(_1654_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(net187),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[5] ),
    .S(_1595_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _3349_ (.A(_1655_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _3350_ (.A0(net181),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[6] ),
    .S(_1595_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _3351_ (.A(_1656_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _3352_ (.A0(net175),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[7] ),
    .S(_1595_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _3353_ (.A(_1657_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _3354_ (.A0(net169),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[8] ),
    .S(_1595_),
    .X(_1658_));
 sky130_fd_sc_hd__clkbuf_1 _3355_ (.A(_1658_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _3356_ (.A0(net164),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[9] ),
    .S(_0422_),
    .X(_1659_));
 sky130_fd_sc_hd__clkbuf_1 _3357_ (.A(_1659_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(\cpu.ALU_OUT_MEMORY_4[10] ),
    .A1(\cpu.REG_WRITE_DATA_WRITEBACK_5[10] ),
    .S(_0422_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3359_ (.A(_1660_),
    .X(_0162_));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.CLK(clknet_leaf_32_CLK),
    .D(_0029_),
    .Q(\cpu.INSTRUCTION_DECODE_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.CLK(clknet_leaf_42_CLK),
    .D(_0030_),
    .Q(\cpu.INSTRUCTION_DECODE_2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.CLK(clknet_leaf_41_CLK),
    .D(_0031_),
    .Q(\cpu.INSTRUCTION_DECODE_2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.CLK(clknet_leaf_33_CLK),
    .D(_0032_),
    .Q(\cpu.INSTRUCTION_DECODE_2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.CLK(clknet_leaf_33_CLK),
    .D(_0033_),
    .Q(\cpu.INSTRUCTION_DECODE_2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.CLK(clknet_leaf_32_CLK),
    .D(_0034_),
    .Q(\cpu.INSTRUCTION_DECODE_2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.CLK(clknet_leaf_0_CLK),
    .D(_0035_),
    .Q(\cpu.INSTRUCTION_DECODE_2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.CLK(clknet_leaf_42_CLK),
    .D(_0036_),
    .Q(\cpu.INSTRUCTION_DECODE_2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.CLK(clknet_leaf_2_CLK),
    .D(_0037_),
    .Q(\cpu.INSTRUCTION_DECODE_2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.CLK(clknet_leaf_33_CLK),
    .D(_0038_),
    .Q(\cpu.INSTRUCTION_DECODE_2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.CLK(clknet_leaf_34_CLK),
    .D(_0039_),
    .Q(\cpu.INSTRUCTION_DECODE_2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3371_ (.CLK(clknet_leaf_32_CLK),
    .D(_0040_),
    .Q(\cpu.R1_PIPELINE[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3372_ (.CLK(clknet_leaf_41_CLK),
    .D(_0041_),
    .Q(\cpu.INSTRUCTION_DECODE_2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3373_ (.CLK(clknet_leaf_33_CLK),
    .D(_0005_),
    .Q(\cpu.TYPE_PIPELINE[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3374_ (.CLK(clknet_leaf_35_CLK),
    .D(_0006_),
    .Q(\cpu.TYPE_PIPELINE[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3375_ (.CLK(clknet_leaf_35_CLK),
    .D(_0007_),
    .Q(\cpu.TYPE_PIPELINE[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.CLK(clknet_leaf_33_CLK),
    .D(_0008_),
    .Q(\cpu.TYPE_PIPELINE[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.CLK(clknet_leaf_33_CLK),
    .D(_0009_),
    .Q(\cpu.TYPE_PIPELINE[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.CLK(clknet_leaf_42_CLK),
    .D(_0000_),
    .Q(\cpu.TYPE_PIPELINE[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.CLK(clknet_leaf_43_CLK),
    .D(net253),
    .Q(\cpu.TYPE_PIPELINE[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3380_ (.CLK(clknet_leaf_42_CLK),
    .D(_0002_),
    .Q(\cpu.TYPE_PIPELINE[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3381_ (.CLK(clknet_leaf_42_CLK),
    .D(_0003_),
    .Q(\cpu.TYPE_PIPELINE[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.CLK(clknet_leaf_42_CLK),
    .D(_0004_),
    .Q(\cpu.TYPE_PIPELINE[0][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3383_ (.D(net145),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3384_ (.D(net158),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3385_ (.D(net153),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3386_ (.D(net157),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3387_ (.D(net150),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3388_ (.D(net142),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3389_ (.D(net151),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3390_ (.D(net147),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3391_ (.D(net129),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3392_ (.D(net132),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3393_ (.D(net133),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3394_ (.D(net135),
    .GATE_N(net59),
    .Q(\cpu.regFile.REGISTERS[10][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3395_ (.D(net123),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3396_ (.D(net138),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3397_ (.D(net96),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3398_ (.D(net140),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3399_ (.D(net113),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3400_ (.D(net115),
    .GATE_N(net58),
    .Q(\cpu.regFile.REGISTERS[10][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3401_ (.D(net98),
    .GATE_N(net57),
    .Q(\cpu.regFile.REGISTERS[10][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3402_ (.D(net100),
    .GATE_N(net57),
    .Q(\cpu.regFile.REGISTERS[10][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3403_ (.D(net117),
    .GATE_N(net57),
    .Q(\cpu.regFile.REGISTERS[10][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3404_ (.D(net128),
    .GATE_N(net57),
    .Q(\cpu.regFile.REGISTERS[10][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3405_ (.D(net119),
    .GATE_N(net57),
    .Q(\cpu.regFile.REGISTERS[10][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3406_ (.D(net121),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3407_ (.D(net80),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3408_ (.D(net83),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3409_ (.D(net84),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3410_ (.D(net86),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3411_ (.D(net88),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3412_ (.D(net90),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3413_ (.D(net92),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3414_ (.D(net95),
    .GATE_N(net56),
    .Q(\cpu.regFile.REGISTERS[10][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3415_ (.D(net144),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3416_ (.D(net158),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3417_ (.D(net153),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3418_ (.D(net157),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3419_ (.D(net149),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3420_ (.D(net141),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3421_ (.D(net151),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3422_ (.D(net147),
    .GATE_N(net112),
    .Q(\cpu.regFile.REGISTERS[15][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3423_ (.D(net129),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3424_ (.D(net131),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3425_ (.D(net133),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3426_ (.D(net135),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3427_ (.D(net123),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3428_ (.D(net138),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3429_ (.D(net97),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3430_ (.D(net140),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3431_ (.D(net114),
    .GATE_N(net110),
    .Q(\cpu.regFile.REGISTERS[15][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3432_ (.D(net116),
    .GATE_N(net111),
    .Q(\cpu.regFile.REGISTERS[15][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3433_ (.D(net99),
    .GATE_N(net111),
    .Q(\cpu.regFile.REGISTERS[15][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3434_ (.D(net101),
    .GATE_N(net111),
    .Q(\cpu.regFile.REGISTERS[15][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3435_ (.D(net118),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3436_ (.D(net127),
    .GATE_N(net111),
    .Q(\cpu.regFile.REGISTERS[15][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3437_ (.D(net120),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3438_ (.D(net122),
    .GATE_N(net111),
    .Q(\cpu.regFile.REGISTERS[15][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3439_ (.D(net81),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3440_ (.D(net83),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3441_ (.D(net85),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3442_ (.D(net87),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3443_ (.D(net89),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3444_ (.D(net91),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3445_ (.D(net93),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3446_ (.D(net95),
    .GATE_N(net109),
    .Q(\cpu.regFile.REGISTERS[15][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3447_ (.D(net144),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3448_ (.D(net158),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3449_ (.D(net153),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3450_ (.D(net156),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3451_ (.D(net150),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3452_ (.D(net142),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3453_ (.D(net151),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3454_ (.D(net148),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3455_ (.D(net129),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3456_ (.D(net132),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3457_ (.D(net133),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3458_ (.D(net135),
    .GATE_N(_0024_),
    .Q(\cpu.regFile.REGISTERS[11][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3459_ (.D(net123),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3460_ (.D(net137),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3461_ (.D(net96),
    .GATE_N(_0024_),
    .Q(\cpu.regFile.REGISTERS[11][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3462_ (.D(net140),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3463_ (.D(net113),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3464_ (.D(net115),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3465_ (.D(net99),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3466_ (.D(net100),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3467_ (.D(net117),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3468_ (.D(net127),
    .GATE_N(net106),
    .Q(\cpu.regFile.REGISTERS[11][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3469_ (.D(net119),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3470_ (.D(net121),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3471_ (.D(net80),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3472_ (.D(net82),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3473_ (.D(net84),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3474_ (.D(net86),
    .GATE_N(net108),
    .Q(\cpu.regFile.REGISTERS[11][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3475_ (.D(net88),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3476_ (.D(net90),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3477_ (.D(net93),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3478_ (.D(net95),
    .GATE_N(net107),
    .Q(\cpu.regFile.REGISTERS[11][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3479_ (.D(net144),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3480_ (.D(net159),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3481_ (.D(net153),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3482_ (.D(net156),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3483_ (.D(net149),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3484_ (.D(net141),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3485_ (.D(net151),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3486_ (.D(net148),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3487_ (.D(net129),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3488_ (.D(net131),
    .GATE_N(net55),
    .Q(\cpu.regFile.REGISTERS[12][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3489_ (.D(net134),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3490_ (.D(net136),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3491_ (.D(net124),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3492_ (.D(net137),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3493_ (.D(net97),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3494_ (.D(net139),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3495_ (.D(net114),
    .GATE_N(net53),
    .Q(\cpu.regFile.REGISTERS[12][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3496_ (.D(net115),
    .GATE_N(net54),
    .Q(\cpu.regFile.REGISTERS[12][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3497_ (.D(net98),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3498_ (.D(net100),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3499_ (.D(net117),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3500_ (.D(net128),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3501_ (.D(net119),
    .GATE_N(net53),
    .Q(\cpu.regFile.REGISTERS[12][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3502_ (.D(net121),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3503_ (.D(net80),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3504_ (.D(net82),
    .GATE_N(net53),
    .Q(\cpu.regFile.REGISTERS[12][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3505_ (.D(net84),
    .GATE_N(net53),
    .Q(\cpu.regFile.REGISTERS[12][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3506_ (.D(net86),
    .GATE_N(net53),
    .Q(\cpu.regFile.REGISTERS[12][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3507_ (.D(net88),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3508_ (.D(net90),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3509_ (.D(net93),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3510_ (.D(net94),
    .GATE_N(net52),
    .Q(\cpu.regFile.REGISTERS[12][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3511_ (.D(net146),
    .GATE_N(net255),
    .Q(\cpu.regFile.REGISTERS[0][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3512_ (.D(net160),
    .GATE_N(net256),
    .Q(\cpu.regFile.REGISTERS[0][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3513_ (.D(net153),
    .GATE_N(net257),
    .Q(\cpu.regFile.REGISTERS[0][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3514_ (.D(net156),
    .GATE_N(net258),
    .Q(\cpu.regFile.REGISTERS[0][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3515_ (.D(net150),
    .GATE_N(net259),
    .Q(\cpu.regFile.REGISTERS[0][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3516_ (.D(net143),
    .GATE_N(net260),
    .Q(\cpu.regFile.REGISTERS[0][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3517_ (.D(net152),
    .GATE_N(net261),
    .Q(\cpu.regFile.REGISTERS[0][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3518_ (.D(net148),
    .GATE_N(net262),
    .Q(\cpu.regFile.REGISTERS[0][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3519_ (.D(net130),
    .GATE_N(net263),
    .Q(\cpu.regFile.REGISTERS[0][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3520_ (.D(net132),
    .GATE_N(net264),
    .Q(\cpu.regFile.REGISTERS[0][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3521_ (.D(\cpu.REG_WRITE_DATA[10] ),
    .GATE_N(net265),
    .Q(\cpu.regFile.REGISTERS[0][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3522_ (.D(net135),
    .GATE_N(net266),
    .Q(\cpu.regFile.REGISTERS[0][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3523_ (.D(net124),
    .GATE_N(net267),
    .Q(\cpu.regFile.REGISTERS[0][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3524_ (.D(net138),
    .GATE_N(net268),
    .Q(\cpu.regFile.REGISTERS[0][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3525_ (.D(net97),
    .GATE_N(net269),
    .Q(\cpu.regFile.REGISTERS[0][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3526_ (.D(net140),
    .GATE_N(net270),
    .Q(\cpu.regFile.REGISTERS[0][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3527_ (.D(net113),
    .GATE_N(net271),
    .Q(\cpu.regFile.REGISTERS[0][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3528_ (.D(net115),
    .GATE_N(net272),
    .Q(\cpu.regFile.REGISTERS[0][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3529_ (.D(net99),
    .GATE_N(net273),
    .Q(\cpu.regFile.REGISTERS[0][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3530_ (.D(net101),
    .GATE_N(net274),
    .Q(\cpu.regFile.REGISTERS[0][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3531_ (.D(net117),
    .GATE_N(net275),
    .Q(\cpu.regFile.REGISTERS[0][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3532_ (.D(net128),
    .GATE_N(net276),
    .Q(\cpu.regFile.REGISTERS[0][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3533_ (.D(net119),
    .GATE_N(net277),
    .Q(\cpu.regFile.REGISTERS[0][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3534_ (.D(net121),
    .GATE_N(net278),
    .Q(\cpu.regFile.REGISTERS[0][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3535_ (.D(net80),
    .GATE_N(net279),
    .Q(\cpu.regFile.REGISTERS[0][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3536_ (.D(net82),
    .GATE_N(net280),
    .Q(\cpu.regFile.REGISTERS[0][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3537_ (.D(net84),
    .GATE_N(net281),
    .Q(\cpu.regFile.REGISTERS[0][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3538_ (.D(net86),
    .GATE_N(net282),
    .Q(\cpu.regFile.REGISTERS[0][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3539_ (.D(net88),
    .GATE_N(net283),
    .Q(\cpu.regFile.REGISTERS[0][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3540_ (.D(net90),
    .GATE_N(net284),
    .Q(\cpu.regFile.REGISTERS[0][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3541_ (.D(net93),
    .GATE_N(net285),
    .Q(\cpu.regFile.REGISTERS[0][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3542_ (.D(net95),
    .GATE_N(net286),
    .Q(\cpu.regFile.REGISTERS[0][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3543_ (.D(net144),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3544_ (.D(net159),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3545_ (.D(net154),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3546_ (.D(net156),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3547_ (.D(net150),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3548_ (.D(net142),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3549_ (.D(net151),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3550_ (.D(net147),
    .GATE_N(net75),
    .Q(\cpu.regFile.REGISTERS[1][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3551_ (.D(net129),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3552_ (.D(net131),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3553_ (.D(net134),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3554_ (.D(net136),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3555_ (.D(net123),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3556_ (.D(net137),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3557_ (.D(net96),
    .GATE_N(net73),
    .Q(\cpu.regFile.REGISTERS[1][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3558_ (.D(net139),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3559_ (.D(net114),
    .GATE_N(net73),
    .Q(\cpu.regFile.REGISTERS[1][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3560_ (.D(net116),
    .GATE_N(net74),
    .Q(\cpu.regFile.REGISTERS[1][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3561_ (.D(net98),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3562_ (.D(net100),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3563_ (.D(net118),
    .GATE_N(net73),
    .Q(\cpu.regFile.REGISTERS[1][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3564_ (.D(net127),
    .GATE_N(net73),
    .Q(\cpu.regFile.REGISTERS[1][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3565_ (.D(net120),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3566_ (.D(net122),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3567_ (.D(net81),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3568_ (.D(net83),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3569_ (.D(net85),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3570_ (.D(net87),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3571_ (.D(net89),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3572_ (.D(net91),
    .GATE_N(net72),
    .Q(\cpu.regFile.REGISTERS[1][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3573_ (.D(net92),
    .GATE_N(net73),
    .Q(\cpu.regFile.REGISTERS[1][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3574_ (.D(net94),
    .GATE_N(net73),
    .Q(\cpu.regFile.REGISTERS[1][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3575_ (.D(net145),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3576_ (.D(net159),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3577_ (.D(net154),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3578_ (.D(net157),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3579_ (.D(net149),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3580_ (.D(net141),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3581_ (.D(net152),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3582_ (.D(net147),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3583_ (.D(net130),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3584_ (.D(net132),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3585_ (.D(net133),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3586_ (.D(net135),
    .GATE_N(net78),
    .Q(\cpu.regFile.REGISTERS[13][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3587_ (.D(net123),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3588_ (.D(net138),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3589_ (.D(net97),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3590_ (.D(net139),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3591_ (.D(net113),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3592_ (.D(net116),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3593_ (.D(net98),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3594_ (.D(net100),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3595_ (.D(net117),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3596_ (.D(net127),
    .GATE_N(net77),
    .Q(\cpu.regFile.REGISTERS[13][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3597_ (.D(net119),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3598_ (.D(net121),
    .GATE_N(net79),
    .Q(\cpu.regFile.REGISTERS[13][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3599_ (.D(net80),
    .GATE_N(net79),
    .Q(\cpu.regFile.REGISTERS[13][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3600_ (.D(net82),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3601_ (.D(net84),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3602_ (.D(net86),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3603_ (.D(net88),
    .GATE_N(net79),
    .Q(\cpu.regFile.REGISTERS[13][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3604_ (.D(net90),
    .GATE_N(net79),
    .Q(\cpu.regFile.REGISTERS[13][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3605_ (.D(net93),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3606_ (.D(net94),
    .GATE_N(net76),
    .Q(\cpu.regFile.REGISTERS[13][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3607_ (.D(net144),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3608_ (.D(net158),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3609_ (.D(net153),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3610_ (.D(net156),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3611_ (.D(net149),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3612_ (.D(net141),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3613_ (.D(net151),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3614_ (.D(net147),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3615_ (.D(net129),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3616_ (.D(net131),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3617_ (.D(net133),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3618_ (.D(net136),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3619_ (.D(net123),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3620_ (.D(net137),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3621_ (.D(net96),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3622_ (.D(net139),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3623_ (.D(net114),
    .GATE_N(net49),
    .Q(\cpu.regFile.REGISTERS[2][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3624_ (.D(net116),
    .GATE_N(net51),
    .Q(\cpu.regFile.REGISTERS[2][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3625_ (.D(net98),
    .GATE_N(net49),
    .Q(\cpu.regFile.REGISTERS[2][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3626_ (.D(net100),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3627_ (.D(net118),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3628_ (.D(net128),
    .GATE_N(net50),
    .Q(\cpu.regFile.REGISTERS[2][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3629_ (.D(net120),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3630_ (.D(net122),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3631_ (.D(net81),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3632_ (.D(net83),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3633_ (.D(net85),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3634_ (.D(net87),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3635_ (.D(net89),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3636_ (.D(net91),
    .GATE_N(net48),
    .Q(\cpu.regFile.REGISTERS[2][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3637_ (.D(net92),
    .GATE_N(net49),
    .Q(\cpu.regFile.REGISTERS[2][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3638_ (.D(net95),
    .GATE_N(net49),
    .Q(\cpu.regFile.REGISTERS[2][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3639_ (.D(net145),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3640_ (.D(net158),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3641_ (.D(net153),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3642_ (.D(net157),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3643_ (.D(net149),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3644_ (.D(net141),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3645_ (.D(net151),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3646_ (.D(net147),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3647_ (.D(net129),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3648_ (.D(net131),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3649_ (.D(net133),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3650_ (.D(net136),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3651_ (.D(net123),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3652_ (.D(net137),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3653_ (.D(net96),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3654_ (.D(net139),
    .GATE_N(net70),
    .Q(\cpu.regFile.REGISTERS[3][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3655_ (.D(net114),
    .GATE_N(net69),
    .Q(\cpu.regFile.REGISTERS[3][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3656_ (.D(net116),
    .GATE_N(net71),
    .Q(\cpu.regFile.REGISTERS[3][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3657_ (.D(net98),
    .GATE_N(net69),
    .Q(\cpu.regFile.REGISTERS[3][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3658_ (.D(net100),
    .GATE_N(net69),
    .Q(\cpu.regFile.REGISTERS[3][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3659_ (.D(net117),
    .GATE_N(net69),
    .Q(\cpu.regFile.REGISTERS[3][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3660_ (.D(net127),
    .GATE_N(net69),
    .Q(\cpu.regFile.REGISTERS[3][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3661_ (.D(net120),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3662_ (.D(net122),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3663_ (.D(net81),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3664_ (.D(net83),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3665_ (.D(net85),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3666_ (.D(net87),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3667_ (.D(net89),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3668_ (.D(net91),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3669_ (.D(net92),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3670_ (.D(net94),
    .GATE_N(net68),
    .Q(\cpu.regFile.REGISTERS[3][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3671_ (.D(net145),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3672_ (.D(net159),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3673_ (.D(net154),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3674_ (.D(net157),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3675_ (.D(net149),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3676_ (.D(net141),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3677_ (.D(net152),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3678_ (.D(net148),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3679_ (.D(net129),
    .GATE_N(net47),
    .Q(\cpu.regFile.REGISTERS[4][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3680_ (.D(net131),
    .GATE_N(net47),
    .Q(\cpu.regFile.REGISTERS[4][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3681_ (.D(net134),
    .GATE_N(net47),
    .Q(\cpu.regFile.REGISTERS[4][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3682_ (.D(net135),
    .GATE_N(net47),
    .Q(\cpu.regFile.REGISTERS[4][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3683_ (.D(net124),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3684_ (.D(net138),
    .GATE_N(net46),
    .Q(\cpu.regFile.REGISTERS[4][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3685_ (.D(net96),
    .GATE_N(net47),
    .Q(\cpu.regFile.REGISTERS[4][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3686_ (.D(net140),
    .GATE_N(net45),
    .Q(\cpu.regFile.REGISTERS[4][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3687_ (.D(net114),
    .GATE_N(net45),
    .Q(\cpu.regFile.REGISTERS[4][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3688_ (.D(net115),
    .GATE_N(net47),
    .Q(\cpu.regFile.REGISTERS[4][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3689_ (.D(net98),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3690_ (.D(net101),
    .GATE_N(net45),
    .Q(\cpu.regFile.REGISTERS[4][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3691_ (.D(net117),
    .GATE_N(net45),
    .Q(\cpu.regFile.REGISTERS[4][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3692_ (.D(net128),
    .GATE_N(net45),
    .Q(\cpu.regFile.REGISTERS[4][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3693_ (.D(net119),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3694_ (.D(net121),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3695_ (.D(net80),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3696_ (.D(net83),
    .GATE_N(net45),
    .Q(\cpu.regFile.REGISTERS[4][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3697_ (.D(net84),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3698_ (.D(net86),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3699_ (.D(net88),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3700_ (.D(net90),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3701_ (.D(net92),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3702_ (.D(net94),
    .GATE_N(net44),
    .Q(\cpu.regFile.REGISTERS[4][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3703_ (.D(net144),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3704_ (.D(net159),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3705_ (.D(net153),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3706_ (.D(net157),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3707_ (.D(net149),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3708_ (.D(net141),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3709_ (.D(net152),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3710_ (.D(net147),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3711_ (.D(net129),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3712_ (.D(net131),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3713_ (.D(net134),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3714_ (.D(net136),
    .GATE_N(net66),
    .Q(\cpu.regFile.REGISTERS[5][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3715_ (.D(net123),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3716_ (.D(net137),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3717_ (.D(net96),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3718_ (.D(net139),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3719_ (.D(net113),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3720_ (.D(net115),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3721_ (.D(net98),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3722_ (.D(net100),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3723_ (.D(net117),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3724_ (.D(net127),
    .GATE_N(net65),
    .Q(\cpu.regFile.REGISTERS[5][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3725_ (.D(net119),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3726_ (.D(net121),
    .GATE_N(net67),
    .Q(\cpu.regFile.REGISTERS[5][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3727_ (.D(net80),
    .GATE_N(net67),
    .Q(\cpu.regFile.REGISTERS[5][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3728_ (.D(net82),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3729_ (.D(net84),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3730_ (.D(net86),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3731_ (.D(net88),
    .GATE_N(net67),
    .Q(\cpu.regFile.REGISTERS[5][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3732_ (.D(net90),
    .GATE_N(net67),
    .Q(\cpu.regFile.REGISTERS[5][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3733_ (.D(net93),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3734_ (.D(net94),
    .GATE_N(net64),
    .Q(\cpu.regFile.REGISTERS[5][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3735_ (.D(net146),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3736_ (.D(net158),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3737_ (.D(net155),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3738_ (.D(net156),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3739_ (.D(net150),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3740_ (.D(net143),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3741_ (.D(net152),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3742_ (.D(net148),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3743_ (.D(net130),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3744_ (.D(net132),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3745_ (.D(net134),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3746_ (.D(net135),
    .GATE_N(net40),
    .Q(\cpu.regFile.REGISTERS[6][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3747_ (.D(net124),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3748_ (.D(net138),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3749_ (.D(net97),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3750_ (.D(net140),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3751_ (.D(net113),
    .GATE_N(net38),
    .Q(\cpu.regFile.REGISTERS[6][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3752_ (.D(net115),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3753_ (.D(net99),
    .GATE_N(net38),
    .Q(\cpu.regFile.REGISTERS[6][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3754_ (.D(net101),
    .GATE_N(net38),
    .Q(\cpu.regFile.REGISTERS[6][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3755_ (.D(net117),
    .GATE_N(net38),
    .Q(\cpu.regFile.REGISTERS[6][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3756_ (.D(net128),
    .GATE_N(net39),
    .Q(\cpu.regFile.REGISTERS[6][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3757_ (.D(net119),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3758_ (.D(net121),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3759_ (.D(net80),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3760_ (.D(net82),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3761_ (.D(net84),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3762_ (.D(net86),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3763_ (.D(net88),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3764_ (.D(net90),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3765_ (.D(net92),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3766_ (.D(net95),
    .GATE_N(net37),
    .Q(\cpu.regFile.REGISTERS[6][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3767_ (.D(net144),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3768_ (.D(net158),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3769_ (.D(net153),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3770_ (.D(net156),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3771_ (.D(net149),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3772_ (.D(net141),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3773_ (.D(net151),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3774_ (.D(net147),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3775_ (.D(net130),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3776_ (.D(net131),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3777_ (.D(net133),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3778_ (.D(net136),
    .GATE_N(_0027_),
    .Q(\cpu.regFile.REGISTERS[14][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3779_ (.D(net124),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3780_ (.D(net137),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3781_ (.D(net97),
    .GATE_N(_0027_),
    .Q(\cpu.regFile.REGISTERS[14][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3782_ (.D(net139),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3783_ (.D(net113),
    .GATE_N(net43),
    .Q(\cpu.regFile.REGISTERS[14][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3784_ (.D(net116),
    .GATE_N(_0027_),
    .Q(\cpu.regFile.REGISTERS[14][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3785_ (.D(net99),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3786_ (.D(net101),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3787_ (.D(net118),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3788_ (.D(net127),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3789_ (.D(net120),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3790_ (.D(net122),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3791_ (.D(net81),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3792_ (.D(net82),
    .GATE_N(net42),
    .Q(\cpu.regFile.REGISTERS[14][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3793_ (.D(net85),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3794_ (.D(net87),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3795_ (.D(net89),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3796_ (.D(net91),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3797_ (.D(net92),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3798_ (.D(net94),
    .GATE_N(net41),
    .Q(\cpu.regFile.REGISTERS[14][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3799_ (.D(net144),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3800_ (.D(net158),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3801_ (.D(net155),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3802_ (.D(net156),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3803_ (.D(net150),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3804_ (.D(net142),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3805_ (.D(net151),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3806_ (.D(net147),
    .GATE_N(net105),
    .Q(\cpu.regFile.REGISTERS[7][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3807_ (.D(net129),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3808_ (.D(net132),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3809_ (.D(net133),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3810_ (.D(net135),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3811_ (.D(net123),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3812_ (.D(net137),
    .GATE_N(net104),
    .Q(\cpu.regFile.REGISTERS[7][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3813_ (.D(net96),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3814_ (.D(net139),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3815_ (.D(net113),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3816_ (.D(net115),
    .GATE_N(net103),
    .Q(\cpu.regFile.REGISTERS[7][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3817_ (.D(net98),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3818_ (.D(net100),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3819_ (.D(net118),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3820_ (.D(net127),
    .GATE_N(net104),
    .Q(\cpu.regFile.REGISTERS[7][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3821_ (.D(net120),
    .GATE_N(net104),
    .Q(\cpu.regFile.REGISTERS[7][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3822_ (.D(net122),
    .GATE_N(net104),
    .Q(\cpu.regFile.REGISTERS[7][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3823_ (.D(net81),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3824_ (.D(net82),
    .GATE_N(net104),
    .Q(\cpu.regFile.REGISTERS[7][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3825_ (.D(net85),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3826_ (.D(net87),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3827_ (.D(net89),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3828_ (.D(net91),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3829_ (.D(net92),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3830_ (.D(net94),
    .GATE_N(net102),
    .Q(\cpu.regFile.REGISTERS[7][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3831_ (.D(net144),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3832_ (.D(net158),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3833_ (.D(net153),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3834_ (.D(net156),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3835_ (.D(net149),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3836_ (.D(net141),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3837_ (.D(net151),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3838_ (.D(net148),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3839_ (.D(net130),
    .GATE_N(net36),
    .Q(\cpu.regFile.REGISTERS[8][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3840_ (.D(net131),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3841_ (.D(net133),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3842_ (.D(net135),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3843_ (.D(net124),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3844_ (.D(net137),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3845_ (.D(net96),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3846_ (.D(net139),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3847_ (.D(net113),
    .GATE_N(net34),
    .Q(\cpu.regFile.REGISTERS[8][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3848_ (.D(net116),
    .GATE_N(net35),
    .Q(\cpu.regFile.REGISTERS[8][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3849_ (.D(net98),
    .GATE_N(net34),
    .Q(\cpu.regFile.REGISTERS[8][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3850_ (.D(net101),
    .GATE_N(net34),
    .Q(\cpu.regFile.REGISTERS[8][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3851_ (.D(net118),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3852_ (.D(net127),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3853_ (.D(net120),
    .GATE_N(net34),
    .Q(\cpu.regFile.REGISTERS[8][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3854_ (.D(net121),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3855_ (.D(net80),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3856_ (.D(net83),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3857_ (.D(net84),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3858_ (.D(net86),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3859_ (.D(net88),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3860_ (.D(net91),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3861_ (.D(net92),
    .GATE_N(net33),
    .Q(\cpu.regFile.REGISTERS[8][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3862_ (.D(net94),
    .GATE_N(net34),
    .Q(\cpu.regFile.REGISTERS[8][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3863_ (.D(net144),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][0] ));
 sky130_fd_sc_hd__dlxtn_1 _3864_ (.D(net158),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][1] ));
 sky130_fd_sc_hd__dlxtn_1 _3865_ (.D(net154),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][2] ));
 sky130_fd_sc_hd__dlxtn_1 _3866_ (.D(net156),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][3] ));
 sky130_fd_sc_hd__dlxtn_1 _3867_ (.D(net149),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][4] ));
 sky130_fd_sc_hd__dlxtn_1 _3868_ (.D(net141),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][5] ));
 sky130_fd_sc_hd__dlxtn_1 _3869_ (.D(net152),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][6] ));
 sky130_fd_sc_hd__dlxtn_1 _3870_ (.D(net147),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][7] ));
 sky130_fd_sc_hd__dlxtn_1 _3871_ (.D(net130),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][8] ));
 sky130_fd_sc_hd__dlxtn_1 _3872_ (.D(net131),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][9] ));
 sky130_fd_sc_hd__dlxtn_1 _3873_ (.D(net133),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][10] ));
 sky130_fd_sc_hd__dlxtn_1 _3874_ (.D(net135),
    .GATE_N(net63),
    .Q(\cpu.regFile.REGISTERS[9][11] ));
 sky130_fd_sc_hd__dlxtn_1 _3875_ (.D(net123),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][12] ));
 sky130_fd_sc_hd__dlxtn_1 _3876_ (.D(net137),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][13] ));
 sky130_fd_sc_hd__dlxtn_1 _3877_ (.D(net96),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][14] ));
 sky130_fd_sc_hd__dlxtn_1 _3878_ (.D(net139),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][15] ));
 sky130_fd_sc_hd__dlxtn_1 _3879_ (.D(net114),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][16] ));
 sky130_fd_sc_hd__dlxtn_1 _3880_ (.D(net115),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][17] ));
 sky130_fd_sc_hd__dlxtn_1 _3881_ (.D(net99),
    .GATE_N(net61),
    .Q(\cpu.regFile.REGISTERS[9][18] ));
 sky130_fd_sc_hd__dlxtn_1 _3882_ (.D(net100),
    .GATE_N(net61),
    .Q(\cpu.regFile.REGISTERS[9][19] ));
 sky130_fd_sc_hd__dlxtn_1 _3883_ (.D(net118),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][20] ));
 sky130_fd_sc_hd__dlxtn_1 _3884_ (.D(net127),
    .GATE_N(net62),
    .Q(\cpu.regFile.REGISTERS[9][21] ));
 sky130_fd_sc_hd__dlxtn_1 _3885_ (.D(net119),
    .GATE_N(net61),
    .Q(\cpu.regFile.REGISTERS[9][22] ));
 sky130_fd_sc_hd__dlxtn_1 _3886_ (.D(net122),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][23] ));
 sky130_fd_sc_hd__dlxtn_1 _3887_ (.D(net81),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][24] ));
 sky130_fd_sc_hd__dlxtn_1 _3888_ (.D(net82),
    .GATE_N(net61),
    .Q(\cpu.regFile.REGISTERS[9][25] ));
 sky130_fd_sc_hd__dlxtn_1 _3889_ (.D(net85),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][26] ));
 sky130_fd_sc_hd__dlxtn_1 _3890_ (.D(net87),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][27] ));
 sky130_fd_sc_hd__dlxtn_1 _3891_ (.D(net89),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][28] ));
 sky130_fd_sc_hd__dlxtn_1 _3892_ (.D(net90),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][29] ));
 sky130_fd_sc_hd__dlxtn_1 _3893_ (.D(net92),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][30] ));
 sky130_fd_sc_hd__dlxtn_1 _3894_ (.D(net94),
    .GATE_N(net60),
    .Q(\cpu.regFile.REGISTERS[9][31] ));
 sky130_fd_sc_hd__dlxtn_1 _3895_ (.D(_0163_),
    .GATE_N(net221),
    .Q(\cpu.ALU_OUT[0] ));
 sky130_fd_sc_hd__dlxtn_1 _3896_ (.D(_0174_),
    .GATE_N(net222),
    .Q(\cpu.ALU_OUT[1] ));
 sky130_fd_sc_hd__dlxtn_1 _3897_ (.D(_0185_),
    .GATE_N(net223),
    .Q(\cpu.ALU_OUT[2] ));
 sky130_fd_sc_hd__dlxtn_1 _3898_ (.D(_0188_),
    .GATE_N(net224),
    .Q(\cpu.ALU_OUT[3] ));
 sky130_fd_sc_hd__dlxtn_1 _3899_ (.D(_0189_),
    .GATE_N(net225),
    .Q(\cpu.ALU_OUT[4] ));
 sky130_fd_sc_hd__dlxtn_1 _3900_ (.D(_0190_),
    .GATE_N(net226),
    .Q(\cpu.ALU_OUT[5] ));
 sky130_fd_sc_hd__dlxtn_1 _3901_ (.D(_0191_),
    .GATE_N(net227),
    .Q(\cpu.ALU_OUT[6] ));
 sky130_fd_sc_hd__dlxtn_1 _3902_ (.D(_0192_),
    .GATE_N(net228),
    .Q(\cpu.ALU_OUT[7] ));
 sky130_fd_sc_hd__dlxtn_2 _3903_ (.D(_0193_),
    .GATE_N(net229),
    .Q(\cpu.ALU_OUT[8] ));
 sky130_fd_sc_hd__dlxtn_1 _3904_ (.D(_0194_),
    .GATE_N(net230),
    .Q(\cpu.ALU_OUT[9] ));
 sky130_fd_sc_hd__dlxtn_1 _3905_ (.D(_0164_),
    .GATE_N(net231),
    .Q(\cpu.ALU_OUT[10] ));
 sky130_fd_sc_hd__dlxtn_1 _3906_ (.D(_0165_),
    .GATE_N(net232),
    .Q(\cpu.ALU_OUT[11] ));
 sky130_fd_sc_hd__dlxtn_1 _3907_ (.D(_0166_),
    .GATE_N(net233),
    .Q(\cpu.ALU_OUT[12] ));
 sky130_fd_sc_hd__dlxtn_1 _3908_ (.D(_0167_),
    .GATE_N(net234),
    .Q(\cpu.ALU_OUT[13] ));
 sky130_fd_sc_hd__dlxtn_1 _3909_ (.D(_0168_),
    .GATE_N(net235),
    .Q(\cpu.ALU_OUT[14] ));
 sky130_fd_sc_hd__dlxtn_1 _3910_ (.D(_0169_),
    .GATE_N(net236),
    .Q(\cpu.ALU_OUT[15] ));
 sky130_fd_sc_hd__dlxtn_1 _3911_ (.D(_0170_),
    .GATE_N(net237),
    .Q(\cpu.ALU_OUT[16] ));
 sky130_fd_sc_hd__dlxtn_1 _3912_ (.D(_0171_),
    .GATE_N(net238),
    .Q(\cpu.ALU_OUT[17] ));
 sky130_fd_sc_hd__dlxtn_1 _3913_ (.D(_0172_),
    .GATE_N(net239),
    .Q(\cpu.ALU_OUT[18] ));
 sky130_fd_sc_hd__dlxtn_1 _3914_ (.D(_0173_),
    .GATE_N(net240),
    .Q(\cpu.ALU_OUT[19] ));
 sky130_fd_sc_hd__dlxtn_1 _3915_ (.D(_0175_),
    .GATE_N(net241),
    .Q(\cpu.ALU_OUT[20] ));
 sky130_fd_sc_hd__dlxtn_1 _3916_ (.D(_0176_),
    .GATE_N(net242),
    .Q(\cpu.ALU_OUT[21] ));
 sky130_fd_sc_hd__dlxtn_1 _3917_ (.D(_0177_),
    .GATE_N(net243),
    .Q(\cpu.ALU_OUT[22] ));
 sky130_fd_sc_hd__dlxtn_1 _3918_ (.D(_0178_),
    .GATE_N(net244),
    .Q(\cpu.ALU_OUT[23] ));
 sky130_fd_sc_hd__dlxtn_1 _3919_ (.D(_0179_),
    .GATE_N(net245),
    .Q(\cpu.ALU_OUT[24] ));
 sky130_fd_sc_hd__dlxtn_1 _3920_ (.D(_0180_),
    .GATE_N(net246),
    .Q(\cpu.ALU_OUT[25] ));
 sky130_fd_sc_hd__dlxtn_1 _3921_ (.D(_0181_),
    .GATE_N(net247),
    .Q(\cpu.ALU_OUT[26] ));
 sky130_fd_sc_hd__dlxtn_1 _3922_ (.D(_0182_),
    .GATE_N(net248),
    .Q(\cpu.ALU_OUT[27] ));
 sky130_fd_sc_hd__dlxtn_1 _3923_ (.D(_0183_),
    .GATE_N(net249),
    .Q(\cpu.ALU_OUT[28] ));
 sky130_fd_sc_hd__dlxtn_1 _3924_ (.D(_0184_),
    .GATE_N(net250),
    .Q(\cpu.ALU_OUT[29] ));
 sky130_fd_sc_hd__dlxtn_1 _3925_ (.D(_0186_),
    .GATE_N(net251),
    .Q(\cpu.ALU_OUT[30] ));
 sky130_fd_sc_hd__dlxtn_1 _3926_ (.D(_0187_),
    .GATE_N(net252),
    .Q(\cpu.ALU_OUT[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3927_ (.CLK(clknet_leaf_31_CLK),
    .D(net293),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3928_ (.CLK(clknet_leaf_30_CLK),
    .D(net288),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3929_ (.CLK(clknet_leaf_30_CLK),
    .D(net291),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3930_ (.CLK(clknet_leaf_28_CLK),
    .D(\cpu.INSTRUCTION_MEMORY_4[11] ),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3931_ (.CLK(clknet_leaf_24_CLK),
    .D(net290),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3932_ (.CLK(clknet_leaf_23_CLK),
    .D(\cpu.INSTRUCTION_MEMORY_4[8] ),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3933_ (.CLK(clknet_leaf_26_CLK),
    .D(net292),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3934_ (.CLK(clknet_leaf_26_CLK),
    .D(net287),
    .Q(\cpu.INSTRUCTION_WRITEBACK_5[10] ));
 sky130_fd_sc_hd__dlxtn_1 _3935_ (.D(_0195_),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[0] ));
 sky130_fd_sc_hd__dlxtn_1 _3936_ (.D(_0202_),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[1] ));
 sky130_fd_sc_hd__dlxtn_1 _3937_ (.D(_0204_),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[2] ));
 sky130_fd_sc_hd__dlxtn_1 _3938_ (.D(_0205_),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[3] ));
 sky130_fd_sc_hd__dlxtn_1 _3939_ (.D(_0206_),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[4] ));
 sky130_fd_sc_hd__dlxtn_1 _3940_ (.D(_0196_),
    .GATE_N(_0012_),
    .Q(\cpu.immediateExtractor.VALUE[11] ));
 sky130_fd_sc_hd__dlxtn_1 _3941_ (.D(_0197_),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[13] ));
 sky130_fd_sc_hd__dlxtn_1 _3942_ (.D(_0198_),
    .GATE_N(net126),
    .Q(\cpu.immediateExtractor.VALUE[16] ));
 sky130_fd_sc_hd__dlxtn_1 _3943_ (.D(_0203_),
    .GATE_N(_0012_),
    .Q(\cpu.immediateExtractor.VALUE[10] ));
 sky130_fd_sc_hd__dlxtn_1 _3944_ (.D(_0199_),
    .GATE_N(net126),
    .Q(\cpu.immediateExtractor.VALUE[20] ));
 sky130_fd_sc_hd__dlxtn_1 _3945_ (.D(_0200_),
    .GATE_N(net126),
    .Q(\cpu.immediateExtractor.VALUE[21] ));
 sky130_fd_sc_hd__dlxtn_1 _3946_ (.D(_0201_),
    .GATE_N(net126),
    .Q(\cpu.immediateExtractor.VALUE[22] ));
 sky130_fd_sc_hd__dlxtn_1 _3947_ (.D(\cpu.INSTRUCTION_EXECUTE_3[11] ),
    .GATE_N(net125),
    .Q(\cpu.immediateExtractor.VALUE[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3948_ (.CLK(clknet_leaf_31_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[0] ),
    .Q(\cpu.INSTRUCTION_MEMORY_4[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3949_ (.CLK(clknet_leaf_29_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[4] ),
    .Q(\cpu.INSTRUCTION_MEMORY_4[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3950_ (.CLK(clknet_leaf_30_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[5] ),
    .Q(\cpu.INSTRUCTION_MEMORY_4[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3951_ (.CLK(clknet_leaf_31_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[11] ),
    .Q(\cpu.INSTRUCTION_MEMORY_4[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3952_ (.CLK(clknet_leaf_25_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[7] ),
    .Q(\cpu.INSTRUCTION_MEMORY_4[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3953_ (.CLK(clknet_leaf_26_CLK),
    .D(net289),
    .Q(\cpu.INSTRUCTION_MEMORY_4[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3954_ (.CLK(clknet_leaf_26_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[9] ),
    .Q(\cpu.INSTRUCTION_MEMORY_4[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3955_ (.CLK(clknet_leaf_28_CLK),
    .D(net294),
    .Q(\cpu.INSTRUCTION_MEMORY_4[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3956_ (.CLK(clknet_leaf_30_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[7] ),
    .Q(\cpu.RD_PIPELINE[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3957_ (.CLK(clknet_leaf_29_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[8] ),
    .Q(\cpu.RD_PIPELINE[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3958_ (.CLK(clknet_leaf_30_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[9] ),
    .Q(\cpu.RD_PIPELINE[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3959_ (.CLK(clknet_leaf_29_CLK),
    .D(net296),
    .Q(\cpu.RD_PIPELINE[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3960_ (.CLK(clknet_leaf_29_CLK),
    .D(\cpu.INSTRUCTION_EXECUTE_3[11] ),
    .Q(\cpu.RD_PIPELINE[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3961_ (.CLK(clknet_leaf_34_CLK),
    .D(_0042_),
    .Q(\cpu.PC_EXECUTE_3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3962_ (.CLK(clknet_leaf_34_CLK),
    .D(_0043_),
    .Q(\cpu.PC_EXECUTE_3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3963_ (.CLK(clknet_leaf_41_CLK),
    .D(_0044_),
    .Q(\cpu.PC_EXECUTE_3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3964_ (.CLK(clknet_leaf_40_CLK),
    .D(_0045_),
    .Q(\cpu.PC_EXECUTE_3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3965_ (.CLK(clknet_leaf_40_CLK),
    .D(_0046_),
    .Q(\cpu.PC_EXECUTE_3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3966_ (.CLK(clknet_leaf_39_CLK),
    .D(_0047_),
    .Q(\cpu.PC_EXECUTE_3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3967_ (.CLK(clknet_leaf_38_CLK),
    .D(_0048_),
    .Q(\cpu.PC_EXECUTE_3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3968_ (.CLK(clknet_leaf_37_CLK),
    .D(_0049_),
    .Q(\cpu.PC_EXECUTE_3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3969_ (.CLK(clknet_leaf_37_CLK),
    .D(_0050_),
    .Q(\cpu.PC_EXECUTE_3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3970_ (.CLK(clknet_leaf_40_CLK),
    .D(_0051_),
    .Q(\cpu.PC_EXECUTE_3[9] ));
 sky130_fd_sc_hd__dfxtp_4 _3971_ (.CLK(clknet_leaf_26_CLK),
    .D(_0052_),
    .Q(net1));
 sky130_fd_sc_hd__dfxtp_4 _3972_ (.CLK(clknet_leaf_42_CLK),
    .D(_0053_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_4 _3973_ (.CLK(clknet_leaf_23_CLK),
    .D(_0054_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_4 _3974_ (.CLK(clknet_leaf_26_CLK),
    .D(_0055_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_4 _3975_ (.CLK(clknet_leaf_0_CLK),
    .D(_0056_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_4 _3976_ (.CLK(clknet_leaf_31_CLK),
    .D(_0057_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _3977_ (.CLK(clknet_leaf_23_CLK),
    .D(_0058_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_4 _3978_ (.CLK(clknet_leaf_0_CLK),
    .D(_0059_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_4 _3979_ (.CLK(clknet_leaf_2_CLK),
    .D(_0060_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_4 _3980_ (.CLK(clknet_leaf_23_CLK),
    .D(_0061_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _3981_ (.CLK(clknet_2_0__leaf_CLK),
    .D(_0062_),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_4 _3982_ (.CLK(clknet_leaf_24_CLK),
    .D(_0063_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_4 _3983_ (.CLK(clknet_leaf_25_CLK),
    .D(_0064_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_2 _3984_ (.CLK(clknet_leaf_7_CLK),
    .D(_0065_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_4 _3985_ (.CLK(clknet_leaf_24_CLK),
    .D(_0066_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_2 _3986_ (.CLK(clknet_leaf_11_CLK),
    .D(_0067_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_4 _3987_ (.CLK(clknet_leaf_7_CLK),
    .D(_0068_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _3988_ (.CLK(clknet_leaf_11_CLK),
    .D(_0069_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_4 _3989_ (.CLK(clknet_leaf_7_CLK),
    .D(_0070_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_4 _3990_ (.CLK(clknet_2_0__leaf_CLK),
    .D(_0071_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_4 _3991_ (.CLK(clknet_leaf_14_CLK),
    .D(_0072_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_4 _3992_ (.CLK(clknet_leaf_14_CLK),
    .D(_0073_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_4 _3993_ (.CLK(clknet_leaf_21_CLK),
    .D(_0074_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_4 _3994_ (.CLK(clknet_leaf_37_CLK),
    .D(_0075_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _3995_ (.CLK(clknet_leaf_15_CLK),
    .D(_0076_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_4 _3996_ (.CLK(clknet_leaf_37_CLK),
    .D(_0077_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_2 _3997_ (.CLK(clknet_leaf_13_CLK),
    .D(_0078_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_4 _3998_ (.CLK(clknet_leaf_37_CLK),
    .D(_0079_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_2 _3999_ (.CLK(clknet_leaf_21_CLK),
    .D(_0080_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_4 _4000_ (.CLK(clknet_leaf_37_CLK),
    .D(_0081_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_2 _4001_ (.CLK(clknet_leaf_21_CLK),
    .D(_0082_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_4 _4002_ (.CLK(clknet_leaf_17_CLK),
    .D(_0083_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _4003_ (.CLK(clknet_leaf_34_CLK),
    .D(_0084_),
    .Q(\cpu.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4004_ (.CLK(clknet_leaf_34_CLK),
    .D(_0085_),
    .Q(\cpu.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4005_ (.CLK(clknet_leaf_26_CLK),
    .D(net290),
    .Q(\cpu.RD_PIPELINE[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4006_ (.CLK(clknet_leaf_26_CLK),
    .D(\cpu.INSTRUCTION_MEMORY_4[8] ),
    .Q(\cpu.RD_PIPELINE[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4007_ (.CLK(clknet_leaf_26_CLK),
    .D(net292),
    .Q(\cpu.RD_PIPELINE[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4008_ (.CLK(clknet_leaf_28_CLK),
    .D(net287),
    .Q(\cpu.RD_PIPELINE[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4009_ (.CLK(clknet_leaf_28_CLK),
    .D(\cpu.INSTRUCTION_MEMORY_4[11] ),
    .Q(\cpu.RD_PIPELINE[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4010_ (.CLK(clknet_leaf_34_CLK),
    .D(\cpu.ALU_OUT[0] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4011_ (.CLK(clknet_leaf_34_CLK),
    .D(\cpu.ALU_OUT[1] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4012_ (.CLK(clknet_leaf_34_CLK),
    .D(\cpu.ALU_OUT[2] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4013_ (.CLK(clknet_leaf_40_CLK),
    .D(\cpu.ALU_OUT[3] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4014_ (.CLK(clknet_leaf_40_CLK),
    .D(\cpu.ALU_OUT[4] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4015_ (.CLK(clknet_leaf_34_CLK),
    .D(\cpu.ALU_OUT[5] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4016_ (.CLK(clknet_leaf_34_CLK),
    .D(\cpu.ALU_OUT[6] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4017_ (.CLK(clknet_leaf_36_CLK),
    .D(\cpu.ALU_OUT[7] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4018_ (.CLK(clknet_leaf_34_CLK),
    .D(\cpu.ALU_OUT[8] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4019_ (.CLK(clknet_leaf_36_CLK),
    .D(\cpu.ALU_OUT[9] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4020_ (.CLK(clknet_leaf_19_CLK),
    .D(\cpu.ALU_OUT[10] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4021_ (.CLK(clknet_leaf_19_CLK),
    .D(\cpu.ALU_OUT[11] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4022_ (.CLK(clknet_leaf_9_CLK),
    .D(\cpu.ALU_OUT[12] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4023_ (.CLK(clknet_leaf_18_CLK),
    .D(\cpu.ALU_OUT[13] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4024_ (.CLK(clknet_leaf_8_CLK),
    .D(\cpu.ALU_OUT[14] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4025_ (.CLK(clknet_leaf_18_CLK),
    .D(\cpu.ALU_OUT[15] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4026_ (.CLK(clknet_leaf_17_CLK),
    .D(\cpu.ALU_OUT[16] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4027_ (.CLK(clknet_leaf_9_CLK),
    .D(\cpu.ALU_OUT[17] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4028_ (.CLK(clknet_leaf_18_CLK),
    .D(\cpu.ALU_OUT[18] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4029_ (.CLK(clknet_leaf_17_CLK),
    .D(\cpu.ALU_OUT[19] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4030_ (.CLK(clknet_leaf_17_CLK),
    .D(\cpu.ALU_OUT[20] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4031_ (.CLK(clknet_leaf_17_CLK),
    .D(\cpu.ALU_OUT[21] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4032_ (.CLK(clknet_leaf_17_CLK),
    .D(\cpu.ALU_OUT[22] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4033_ (.CLK(clknet_leaf_16_CLK),
    .D(\cpu.ALU_OUT[23] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4034_ (.CLK(clknet_leaf_16_CLK),
    .D(\cpu.ALU_OUT[24] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4035_ (.CLK(clknet_leaf_15_CLK),
    .D(\cpu.ALU_OUT[25] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4036_ (.CLK(clknet_leaf_15_CLK),
    .D(\cpu.ALU_OUT[26] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4037_ (.CLK(clknet_leaf_15_CLK),
    .D(\cpu.ALU_OUT[27] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4038_ (.CLK(clknet_leaf_15_CLK),
    .D(\cpu.ALU_OUT[28] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4039_ (.CLK(clknet_leaf_16_CLK),
    .D(\cpu.ALU_OUT[29] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4040_ (.CLK(clknet_leaf_15_CLK),
    .D(\cpu.ALU_OUT[30] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4041_ (.CLK(clknet_leaf_15_CLK),
    .D(\cpu.ALU_OUT[31] ),
    .Q(\cpu.ALU_OUT_MEMORY_4[31] ));
 sky130_fd_sc_hd__dfxtp_2 _4042_ (.CLK(clknet_leaf_35_CLK),
    .D(\cpu.PC_EXECUTE_3[0] ),
    .Q(\cpu.PC_MEMORY_4[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4043_ (.CLK(clknet_leaf_35_CLK),
    .D(\cpu.PC_EXECUTE_3[1] ),
    .Q(\cpu.PC_MEMORY_4[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4044_ (.CLK(clknet_leaf_41_CLK),
    .D(\cpu.PC_EXECUTE_3[2] ),
    .Q(\cpu.PC_MEMORY_4[2] ));
 sky130_fd_sc_hd__dfxtp_2 _4045_ (.CLK(clknet_leaf_40_CLK),
    .D(\cpu.PC_EXECUTE_3[3] ),
    .Q(\cpu.PC_MEMORY_4[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4046_ (.CLK(clknet_leaf_40_CLK),
    .D(\cpu.PC_EXECUTE_3[4] ),
    .Q(\cpu.PC_MEMORY_4[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4047_ (.CLK(clknet_leaf_38_CLK),
    .D(\cpu.PC_EXECUTE_3[5] ),
    .Q(\cpu.PC_MEMORY_4[5] ));
 sky130_fd_sc_hd__dfxtp_2 _4048_ (.CLK(clknet_leaf_37_CLK),
    .D(\cpu.PC_EXECUTE_3[6] ),
    .Q(\cpu.PC_MEMORY_4[6] ));
 sky130_fd_sc_hd__dfxtp_2 _4049_ (.CLK(clknet_leaf_37_CLK),
    .D(\cpu.PC_EXECUTE_3[7] ),
    .Q(\cpu.PC_MEMORY_4[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4050_ (.CLK(clknet_leaf_37_CLK),
    .D(\cpu.PC_EXECUTE_3[8] ),
    .Q(\cpu.PC_MEMORY_4[8] ));
 sky130_fd_sc_hd__dfxtp_2 _4051_ (.CLK(clknet_leaf_34_CLK),
    .D(net295),
    .Q(\cpu.PC_MEMORY_4[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4052_ (.CLK(clknet_leaf_0_CLK),
    .D(\cpu.R2_DATA[0] ),
    .Q(\cpu.RAM_WRITE_DATA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4053_ (.CLK(clknet_leaf_43_CLK),
    .D(\cpu.R2_DATA[1] ),
    .Q(\cpu.RAM_WRITE_DATA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4054_ (.CLK(clknet_leaf_2_CLK),
    .D(\cpu.R2_DATA[2] ),
    .Q(\cpu.RAM_WRITE_DATA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4055_ (.CLK(clknet_leaf_2_CLK),
    .D(\cpu.R2_DATA[3] ),
    .Q(\cpu.RAM_WRITE_DATA[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4056_ (.CLK(clknet_leaf_0_CLK),
    .D(\cpu.R2_DATA[4] ),
    .Q(\cpu.RAM_WRITE_DATA[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4057_ (.CLK(clknet_leaf_2_CLK),
    .D(\cpu.R2_DATA[5] ),
    .Q(\cpu.RAM_WRITE_DATA[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4058_ (.CLK(clknet_leaf_31_CLK),
    .D(\cpu.R2_DATA[6] ),
    .Q(\cpu.RAM_WRITE_DATA[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4059_ (.CLK(clknet_leaf_2_CLK),
    .D(\cpu.R2_DATA[7] ),
    .Q(\cpu.RAM_WRITE_DATA[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4060_ (.CLK(clknet_leaf_33_CLK),
    .D(_0086_),
    .Q(\cpu.INSTRUCTION_DECODE_2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4061_ (.CLK(clknet_leaf_8_CLK),
    .D(_0087_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4062_ (.CLK(clknet_leaf_10_CLK),
    .D(_0088_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4063_ (.CLK(clknet_leaf_10_CLK),
    .D(_0089_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4064_ (.CLK(clknet_leaf_9_CLK),
    .D(_0090_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4065_ (.CLK(clknet_leaf_9_CLK),
    .D(_0091_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4066_ (.CLK(clknet_leaf_11_CLK),
    .D(_0092_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4067_ (.CLK(clknet_leaf_9_CLK),
    .D(_0093_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4068_ (.CLK(clknet_leaf_11_CLK),
    .D(_0094_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4069_ (.CLK(clknet_leaf_12_CLK),
    .D(_0095_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4070_ (.CLK(clknet_leaf_12_CLK),
    .D(_0096_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4071_ (.CLK(clknet_leaf_11_CLK),
    .D(_0097_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4072_ (.CLK(clknet_leaf_12_CLK),
    .D(_0098_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4073_ (.CLK(clknet_leaf_12_CLK),
    .D(_0099_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4074_ (.CLK(clknet_leaf_13_CLK),
    .D(_0100_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4075_ (.CLK(clknet_leaf_13_CLK),
    .D(_0101_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4076_ (.CLK(clknet_leaf_13_CLK),
    .D(_0102_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4077_ (.CLK(clknet_leaf_15_CLK),
    .D(_0103_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4078_ (.CLK(clknet_leaf_13_CLK),
    .D(_0104_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4079_ (.CLK(clknet_leaf_13_CLK),
    .D(_0105_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4080_ (.CLK(clknet_leaf_13_CLK),
    .D(_0106_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4081_ (.CLK(clknet_leaf_14_CLK),
    .D(_0107_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4082_ (.CLK(clknet_leaf_34_CLK),
    .D(_0108_),
    .Q(\cpu.PC_DECODE_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4083_ (.CLK(clknet_leaf_34_CLK),
    .D(_0109_),
    .Q(\cpu.PC_DECODE_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4084_ (.CLK(clknet_leaf_41_CLK),
    .D(_0110_),
    .Q(\cpu.PC_DECODE_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4085_ (.CLK(clknet_leaf_40_CLK),
    .D(_0111_),
    .Q(\cpu.PC_DECODE_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4086_ (.CLK(clknet_leaf_39_CLK),
    .D(_0112_),
    .Q(\cpu.PC_DECODE_2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4087_ (.CLK(clknet_leaf_39_CLK),
    .D(_0113_),
    .Q(\cpu.PC_DECODE_2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4088_ (.CLK(clknet_leaf_38_CLK),
    .D(_0114_),
    .Q(\cpu.PC_DECODE_2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4089_ (.CLK(clknet_leaf_38_CLK),
    .D(_0115_),
    .Q(\cpu.PC_DECODE_2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4090_ (.CLK(clknet_leaf_38_CLK),
    .D(_0116_),
    .Q(\cpu.PC_DECODE_2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4091_ (.CLK(clknet_leaf_39_CLK),
    .D(_0117_),
    .Q(\cpu.PC_DECODE_2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _4092_ (.CLK(clknet_leaf_31_CLK),
    .D(_0118_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4093_ (.CLK(clknet_leaf_35_CLK),
    .D(_0119_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4094_ (.CLK(clknet_leaf_30_CLK),
    .D(_0120_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4095_ (.CLK(clknet_leaf_31_CLK),
    .D(_0121_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4096_ (.CLK(clknet_leaf_29_CLK),
    .D(_0122_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4097_ (.CLK(clknet_leaf_31_CLK),
    .D(_0123_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4098_ (.CLK(clknet_leaf_35_CLK),
    .D(_0124_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[10] ));
 sky130_fd_sc_hd__dfxtp_2 _4099_ (.CLK(clknet_leaf_35_CLK),
    .D(_0125_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4100_ (.CLK(clknet_leaf_25_CLK),
    .D(_0126_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[16] ));
 sky130_fd_sc_hd__dfxtp_2 _4101_ (.CLK(clknet_leaf_26_CLK),
    .D(_0127_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[20] ));
 sky130_fd_sc_hd__dfxtp_4 _4102_ (.CLK(clknet_leaf_25_CLK),
    .D(_0128_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[21] ));
 sky130_fd_sc_hd__dfxtp_4 _4103_ (.CLK(clknet_leaf_2_CLK),
    .D(_0129_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[22] ));
 sky130_fd_sc_hd__dfxtp_2 _4104_ (.CLK(clknet_leaf_31_CLK),
    .D(_0130_),
    .Q(\cpu.INSTRUCTION_EXECUTE_3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4105_ (.CLK(clknet_leaf_30_CLK),
    .D(_0131_),
    .Q(\cpu.R1_PIPELINE[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4106_ (.CLK(clknet_leaf_34_CLK),
    .D(_0132_),
    .Q(\cpu.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4107_ (.CLK(clknet_leaf_40_CLK),
    .D(_0133_),
    .Q(\cpu.PC[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4108_ (.CLK(clknet_leaf_39_CLK),
    .D(_0134_),
    .Q(\cpu.PC[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4109_ (.CLK(clknet_leaf_39_CLK),
    .D(_0135_),
    .Q(\cpu.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4110_ (.CLK(clknet_leaf_38_CLK),
    .D(_0136_),
    .Q(\cpu.PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4111_ (.CLK(clknet_leaf_38_CLK),
    .D(_0137_),
    .Q(\cpu.PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4112_ (.CLK(clknet_leaf_36_CLK),
    .D(_0138_),
    .Q(\cpu.PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4113_ (.CLK(clknet_leaf_38_CLK),
    .D(_0139_),
    .Q(\cpu.PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4114_ (.CLK(clknet_leaf_32_CLK),
    .D(_0140_),
    .Q(\cpu.RD_PIPELINE[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4115_ (.CLK(clknet_leaf_32_CLK),
    .D(_0141_),
    .Q(\cpu.RD_PIPELINE[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4116_ (.CLK(clknet_leaf_1_CLK),
    .D(_0142_),
    .Q(\cpu.RD_PIPELINE[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4117_ (.CLK(clknet_leaf_32_CLK),
    .D(_0143_),
    .Q(\cpu.RD_PIPELINE[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _4118_ (.CLK(clknet_leaf_2_CLK),
    .D(_0144_),
    .Q(\cpu.R2_PIPELINE[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4119_ (.CLK(clknet_leaf_1_CLK),
    .D(_0145_),
    .Q(\cpu.R2_PIPELINE[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4120_ (.CLK(clknet_leaf_1_CLK),
    .D(_0146_),
    .Q(\cpu.R2_PIPELINE[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4121_ (.CLK(clknet_leaf_2_CLK),
    .D(_0147_),
    .Q(\cpu.R2_PIPELINE[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4122_ (.CLK(clknet_leaf_42_CLK),
    .D(_0148_),
    .Q(\cpu.R2_PIPELINE[0][3] ));
 sky130_fd_sc_hd__dfxtp_4 _4123_ (.CLK(clknet_leaf_3_CLK),
    .D(\RAM_READ_DATA[0] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[0] ));
 sky130_fd_sc_hd__dfxtp_4 _4124_ (.CLK(clknet_leaf_3_CLK),
    .D(\RAM_READ_DATA[1] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[1] ));
 sky130_fd_sc_hd__dfxtp_4 _4125_ (.CLK(clknet_leaf_4_CLK),
    .D(\RAM_READ_DATA[2] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[2] ));
 sky130_fd_sc_hd__dfxtp_4 _4126_ (.CLK(clknet_leaf_4_CLK),
    .D(\RAM_READ_DATA[3] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4127_ (.CLK(clknet_leaf_4_CLK),
    .D(\RAM_READ_DATA[4] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4128_ (.CLK(clknet_leaf_5_CLK),
    .D(\RAM_READ_DATA[5] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4129_ (.CLK(clknet_leaf_5_CLK),
    .D(\RAM_READ_DATA[6] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[6] ));
 sky130_fd_sc_hd__dfxtp_4 _4130_ (.CLK(clknet_leaf_5_CLK),
    .D(\RAM_READ_DATA[7] ),
    .Q(\cpu.RAM_READ_DATA_WRITEBACK_5[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4131_ (.CLK(clknet_leaf_30_CLK),
    .D(_0149_),
    .Q(\cpu.R2_PIPELINE[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _4132_ (.CLK(clknet_leaf_30_CLK),
    .D(_0150_),
    .Q(\cpu.R2_PIPELINE[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4133_ (.CLK(clknet_leaf_31_CLK),
    .D(_0151_),
    .Q(\cpu.R2_PIPELINE[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4134_ (.CLK(clknet_leaf_30_CLK),
    .D(_0152_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4135_ (.CLK(clknet_leaf_28_CLK),
    .D(_0153_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4136_ (.CLK(clknet_leaf_28_CLK),
    .D(_0154_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4137_ (.CLK(clknet_2_0__leaf_CLK),
    .D(_0155_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4138_ (.CLK(clknet_leaf_26_CLK),
    .D(_0156_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4139_ (.CLK(clknet_leaf_24_CLK),
    .D(_0157_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4140_ (.CLK(clknet_leaf_24_CLK),
    .D(_0158_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4141_ (.CLK(clknet_leaf_24_CLK),
    .D(_0159_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4142_ (.CLK(clknet_leaf_10_CLK),
    .D(_0160_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4143_ (.CLK(clknet_leaf_8_CLK),
    .D(_0161_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4144_ (.CLK(clknet_leaf_8_CLK),
    .D(_0162_),
    .Q(\cpu.REG_WRITE_DATA_WRITEBACK_5[10] ));
 sky130_fd_sc_hd__conb_1 _3511__255 (.HI(net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__conb_1 _3379__253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 ram_254 (.HI(net254));
 sky130_sram_1kbyte_1r1w_8x1024_8 ram (.csb0(_0010_),
    .csb1(net254),
    .clk0(clknet_2_2__leaf_CLK),
    .clk1(clknet_2_1__leaf_CLK),
    .addr0({net161,
    net167,
    net173,
    net179,
    net185,
    net191,
    net197,
    net203,
    net209,
    net215}),
    .addr1({net162,
    net168,
    net174,
    net180,
    net186,
    net192,
    net198,
    net205,
    net211,
    net217}),
    .din0({\cpu.RAM_WRITE_DATA[7] ,
    \cpu.RAM_WRITE_DATA[6] ,
    \cpu.RAM_WRITE_DATA[5] ,
    \cpu.RAM_WRITE_DATA[4] ,
    \cpu.RAM_WRITE_DATA[3] ,
    \cpu.RAM_WRITE_DATA[2] ,
    \cpu.RAM_WRITE_DATA[1] ,
    \cpu.RAM_WRITE_DATA[0] }),
    .dout1({\RAM_READ_DATA[7] ,
    \RAM_READ_DATA[6] ,
    \RAM_READ_DATA[5] ,
    \RAM_READ_DATA[4] ,
    \RAM_READ_DATA[3] ,
    \RAM_READ_DATA[2] ,
    \RAM_READ_DATA[1] ,
    \RAM_READ_DATA[0] }));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(GPIO[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(GPIO[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(GPIO[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(GPIO[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(GPIO[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(GPIO[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(GPIO[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(GPIO[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(GPIO[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(GPIO[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(GPIO[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(GPIO[1]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(GPIO[20]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(GPIO[21]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(GPIO[22]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(GPIO[23]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(GPIO[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(GPIO[25]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(GPIO[26]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(GPIO[27]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(GPIO[28]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(GPIO[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(GPIO[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(GPIO[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(GPIO[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(GPIO[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(GPIO[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(GPIO[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(GPIO[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(GPIO[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(GPIO[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(GPIO[9]));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(_0021_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(_0019_),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(_0027_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(_0027_),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(_0017_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(_0017_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(_0017_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net51),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(_0015_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(_0025_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(_0025_),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(_0023_),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout57 (.A(_0023_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(_0023_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(_0022_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(_0022_),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(net67),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(_0018_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(_0016_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(_0014_),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(net79),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(_0026_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(\cpu.REG_WRITE_DATA[24] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(\cpu.REG_WRITE_DATA[24] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(\cpu.REG_WRITE_DATA[25] ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(\cpu.REG_WRITE_DATA[25] ),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(\cpu.REG_WRITE_DATA[26] ),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout85 (.A(\cpu.REG_WRITE_DATA[26] ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(\cpu.REG_WRITE_DATA[27] ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(\cpu.REG_WRITE_DATA[27] ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(\cpu.REG_WRITE_DATA[28] ),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout89 (.A(\cpu.REG_WRITE_DATA[28] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(\cpu.REG_WRITE_DATA[29] ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(\cpu.REG_WRITE_DATA[29] ),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(\cpu.REG_WRITE_DATA[30] ),
    .X(net93));
 sky130_fd_sc_hd__buf_2 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(\cpu.REG_WRITE_DATA[31] ),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(\cpu.REG_WRITE_DATA[14] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(\cpu.REG_WRITE_DATA[18] ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 fanout101 (.A(\cpu.REG_WRITE_DATA[19] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(_0020_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(_0024_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(_0024_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(_0024_),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net111),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(_0028_),
    .X(net112));
 sky130_fd_sc_hd__buf_2 fanout113 (.A(\cpu.REG_WRITE_DATA[16] ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(\cpu.REG_WRITE_DATA[16] ),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(\cpu.REG_WRITE_DATA[17] ),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(\cpu.REG_WRITE_DATA[17] ),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(\cpu.REG_WRITE_DATA[20] ),
    .X(net117));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout118 (.A(\cpu.REG_WRITE_DATA[20] ),
    .X(net118));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(\cpu.REG_WRITE_DATA[22] ),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(\cpu.REG_WRITE_DATA[22] ),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(\cpu.REG_WRITE_DATA[23] ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(\cpu.REG_WRITE_DATA[23] ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_2 fanout124 (.A(\cpu.REG_WRITE_DATA[12] ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(_0012_),
    .X(net126));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_2 fanout128 (.A(\cpu.REG_WRITE_DATA[21] ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(\cpu.REG_WRITE_DATA[8] ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(\cpu.REG_WRITE_DATA[9] ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(\cpu.REG_WRITE_DATA[10] ),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(\cpu.REG_WRITE_DATA[11] ),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout136 (.A(\cpu.REG_WRITE_DATA[11] ),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(\cpu.REG_WRITE_DATA[13] ),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(\cpu.REG_WRITE_DATA[15] ),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(\cpu.REG_WRITE_DATA[5] ),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(\cpu.REG_WRITE_DATA[0] ),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(\cpu.REG_WRITE_DATA[7] ),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 fanout150 (.A(\cpu.REG_WRITE_DATA[4] ),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(\cpu.REG_WRITE_DATA[6] ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(\cpu.REG_WRITE_DATA[2] ),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(\cpu.REG_WRITE_DATA[3] ),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout157 (.A(\cpu.REG_WRITE_DATA[3] ),
    .X(net157));
 sky130_fd_sc_hd__buf_2 fanout158 (.A(net160),
    .X(net158));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(\cpu.REG_WRITE_DATA[1] ),
    .X(net160));
 sky130_fd_sc_hd__buf_4 wire161 (.A(net166),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 wire162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 wire163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 wire165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_4 wire166 (.A(\cpu.ALU_OUT_MEMORY_4[9] ),
    .X(net166));
 sky130_fd_sc_hd__buf_4 wire167 (.A(net172),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 wire168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 wire169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 wire171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_4 wire172 (.A(\cpu.ALU_OUT_MEMORY_4[8] ),
    .X(net172));
 sky130_fd_sc_hd__buf_4 wire173 (.A(net178),
    .X(net173));
 sky130_fd_sc_hd__buf_2 wire174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_2 wire175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_4 wire178 (.A(\cpu.ALU_OUT_MEMORY_4[7] ),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 wire179 (.A(net184),
    .X(net179));
 sky130_fd_sc_hd__buf_2 wire180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_2 wire181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 wire182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_4 wire184 (.A(\cpu.ALU_OUT_MEMORY_4[6] ),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 wire185 (.A(net190),
    .X(net185));
 sky130_fd_sc_hd__buf_2 wire186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_2 wire187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 wire188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_4 wire190 (.A(\cpu.ALU_OUT_MEMORY_4[5] ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 wire191 (.A(net196),
    .X(net191));
 sky130_fd_sc_hd__buf_2 wire192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 wire193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_4 wire196 (.A(\cpu.ALU_OUT_MEMORY_4[4] ),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 wire197 (.A(net202),
    .X(net197));
 sky130_fd_sc_hd__buf_2 wire198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 wire199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 wire202 (.A(\cpu.ALU_OUT_MEMORY_4[3] ),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 wire203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 wire204 (.A(net208),
    .X(net204));
 sky130_fd_sc_hd__buf_4 wire205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_4 wire206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 wire207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 wire208 (.A(\cpu.ALU_OUT_MEMORY_4[2] ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 wire209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 wire210 (.A(net214),
    .X(net210));
 sky130_fd_sc_hd__buf_4 wire211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 wire212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 load_slew213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire214 (.A(\cpu.ALU_OUT_MEMORY_4[1] ),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 wire215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 wire216 (.A(net220),
    .X(net216));
 sky130_fd_sc_hd__buf_4 wire217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_4 wire218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 wire219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 wire220 (.A(\cpu.ALU_OUT_MEMORY_4[0] ),
    .X(net220));
 sky130_fd_sc_hd__conb_1 _3895__221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _3896__222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _3897__223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _3898__224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _3899__225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 _3900__226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 _3901__227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 _3902__228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 _3903__229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 _3904__230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 _3905__231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 _3906__232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 _3907__233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 _3908__234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 _3909__235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 _3910__236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 _3911__237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 _3912__238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 _3913__239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 _3914__240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 _3915__241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 _3916__242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 _3917__243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 _3918__244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 _3919__245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 _3920__246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 _3921__247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 _3922__248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 _3923__249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 _3924__250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 _3925__251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 _3926__252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 _3512__256 (.HI(net256));
 sky130_fd_sc_hd__conb_1 _3513__257 (.HI(net257));
 sky130_fd_sc_hd__conb_1 _3514__258 (.HI(net258));
 sky130_fd_sc_hd__conb_1 _3515__259 (.HI(net259));
 sky130_fd_sc_hd__conb_1 _3516__260 (.HI(net260));
 sky130_fd_sc_hd__conb_1 _3517__261 (.HI(net261));
 sky130_fd_sc_hd__conb_1 _3518__262 (.HI(net262));
 sky130_fd_sc_hd__conb_1 _3519__263 (.HI(net263));
 sky130_fd_sc_hd__conb_1 _3520__264 (.HI(net264));
 sky130_fd_sc_hd__conb_1 _3521__265 (.HI(net265));
 sky130_fd_sc_hd__conb_1 _3522__266 (.HI(net266));
 sky130_fd_sc_hd__conb_1 _3523__267 (.HI(net267));
 sky130_fd_sc_hd__conb_1 _3524__268 (.HI(net268));
 sky130_fd_sc_hd__conb_1 _3525__269 (.HI(net269));
 sky130_fd_sc_hd__conb_1 _3526__270 (.HI(net270));
 sky130_fd_sc_hd__conb_1 _3527__271 (.HI(net271));
 sky130_fd_sc_hd__conb_1 _3528__272 (.HI(net272));
 sky130_fd_sc_hd__conb_1 _3529__273 (.HI(net273));
 sky130_fd_sc_hd__conb_1 _3530__274 (.HI(net274));
 sky130_fd_sc_hd__conb_1 _3531__275 (.HI(net275));
 sky130_fd_sc_hd__conb_1 _3532__276 (.HI(net276));
 sky130_fd_sc_hd__conb_1 _3533__277 (.HI(net277));
 sky130_fd_sc_hd__conb_1 _3534__278 (.HI(net278));
 sky130_fd_sc_hd__conb_1 _3535__279 (.HI(net279));
 sky130_fd_sc_hd__conb_1 _3536__280 (.HI(net280));
 sky130_fd_sc_hd__conb_1 _3537__281 (.HI(net281));
 sky130_fd_sc_hd__conb_1 _3538__282 (.HI(net282));
 sky130_fd_sc_hd__conb_1 _3539__283 (.HI(net283));
 sky130_fd_sc_hd__conb_1 _3540__284 (.HI(net284));
 sky130_fd_sc_hd__conb_1 _3541__285 (.HI(net285));
 sky130_fd_sc_hd__conb_1 _3542__286 (.HI(net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_CLK (.A(clknet_2_1__leaf_CLK),
    .X(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_CLK (.A(clknet_2_0__leaf_CLK),
    .X(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_CLK (.A(clknet_2_2__leaf_CLK),
    .X(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_CLK (.A(clknet_2_3__leaf_CLK),
    .X(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_1__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_2__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_3__leaf_CLK));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\cpu.INSTRUCTION_MEMORY_4[10] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\cpu.INSTRUCTION_MEMORY_4[4] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\cpu.INSTRUCTION_EXECUTE_3[8] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\cpu.INSTRUCTION_MEMORY_4[7] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\cpu.INSTRUCTION_MEMORY_4[5] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\cpu.INSTRUCTION_MEMORY_4[9] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\cpu.INSTRUCTION_MEMORY_4[0] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\cpu.INSTRUCTION_EXECUTE_3[10] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\cpu.PC_EXECUTE_3[9] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\cpu.INSTRUCTION_EXECUTE_3[10] ),
    .X(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(CLK));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0027_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0128_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\cpu.ALU_OUT[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\cpu.ALU_OUT[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\cpu.INSTRUCTION_EXECUTE_3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\cpu.INSTRUCTION_EXECUTE_3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\cpu.R2_DATA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\cpu.R2_DATA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\cpu.R2_DATA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\cpu.R2_DATA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\cpu.R2_PIPELINE[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\cpu.RAM_READ_DATA_WRITEBACK_5[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\cpu.REG_WRITE_DATA[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\cpu.REG_WRITE_DATA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\cpu.REG_WRITE_DATA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\cpu.PC_EXECUTE_3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1542 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1599 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1603 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1616 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1662 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1718 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1751 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1763 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1793 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1816 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1828 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1846 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1869 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1946 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1958 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1961 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1981 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1994 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1326 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1347 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1434 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1442 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1459 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1559 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1615 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1627 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1696 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1723 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1731 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1779 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1802 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1889 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1969 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1977 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1389 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1448 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1580 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1592 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1604 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1634 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1642 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1690 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1750 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1774 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1799 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1914 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1346 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1516 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1865 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1963 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1979 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1452 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1486 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1524 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1560 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1577 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1583 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1587 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1596 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1606 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1643 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1773 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1817 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1831 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1837 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1846 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1849 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1857 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1872 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1900 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1970 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1982 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1392 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1404 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1412 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1559 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1583 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1617 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1665 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1684 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1700 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1792 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1887 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1895 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1920 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1947 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1971 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2003 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2027 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1643 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1668 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1691 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1703 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1764 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1776 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1885 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1915 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1923 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1336 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1609 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1626 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1638 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1722 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1734 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1897 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1392 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1415 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1433 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1587 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1599 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1607 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1829 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1833 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1846 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1975 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1991 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2011 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1556 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1571 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1582 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1621 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1688 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1783 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1795 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1803 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1857 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1865 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1945 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1957 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1965 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1986 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1495 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1524 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1605 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1692 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1727 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1745 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1759 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1767 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1802 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1810 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1818 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1829 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1845 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1849 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1858 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1876 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1892 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1912 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1924 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1948 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1968 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2004 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2035 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2047 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2059 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1443 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1536 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1649 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1676 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1694 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1721 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1727 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1740 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1802 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1833 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1887 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1895 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1929 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1947 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1968 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1980 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1989 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1997 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2008 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2020 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2028 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1454 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1463 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1586 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1598 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1606 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1766 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1919 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1927 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1942 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1407 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1449 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1556 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1576 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1609 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1617 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1628 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1640 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1915 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1927 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1931 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1946 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1970 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1478 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1490 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1540 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1552 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1587 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1637 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1666 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1694 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1722 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1773 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1814 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1826 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1834 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1975 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2007 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2017 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2025 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2040 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2052 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1336 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1397 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1415 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1510 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1518 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1611 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1624 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1634 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1658 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1682 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1698 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1721 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1745 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1761 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1771 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1795 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1803 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1835 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1846 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1858 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1886 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1957 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1963 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1976 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1984 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2016 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2024 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1415 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1423 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1538 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1544 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1591 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1643 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1659 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1914 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1946 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1958 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2040 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2052 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1267 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1555 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1562 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1574 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1609 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1620 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1720 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1732 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1744 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1833 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1839 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1877 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1889 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1907 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1923 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1931 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1947 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1971 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1454 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1544 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1556 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1679 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1701 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1714 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1940 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1578 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1590 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1609 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1621 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1733 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1850 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1862 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1874 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1945 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1964 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1972 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1989 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2001 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2007 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2020 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2028 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2125 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1584 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1590 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1596 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1600 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1604 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1637 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1645 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1655 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1663 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1749 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1769 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1790 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1812 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1858 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1882 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1894 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1975 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1991 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1999 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2027 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2039 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1522 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1571 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1575 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1583 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1594 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1615 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1691 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1720 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1732 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1744 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1752 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1813 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1835 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1847 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1859 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1887 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1899 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1911 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1923 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2013 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2025 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2029 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1487 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1499 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1605 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1616 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1681 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1919 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1473 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1615 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1627 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1646 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1677 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1721 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1897 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1912 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1947 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1971 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1574 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1586 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1598 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1610 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1639 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1655 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1817 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1829 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1835 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1849 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1861 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1892 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1912 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1924 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2000 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2012 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1393 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1446 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1458 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1516 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1528 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1552 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1564 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1574 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1578 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1672 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1688 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1777 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1795 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1827 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1840 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1852 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1872 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1886 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1945 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1971 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1982 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1989 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1998 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2002 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2014 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2022 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1477 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1556 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1590 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1602 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1608 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1716 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1761 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1802 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1810 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1825 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1967 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1979 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2011 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2015 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2031 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2055 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1392 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1453 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1595 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1605 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1723 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1731 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1741 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1749 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1889 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1901 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1909 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2003 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2027 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1309 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1330 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1376 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1623 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1625 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1633 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1751 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1919 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2037 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2050 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1393 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1616 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1624 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1634 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1640 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1663 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1675 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1687 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1709 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1736 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1752 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1783 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1802 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1821 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1833 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1848 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1864 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1891 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1916 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1928 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1947 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1970 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2059 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2083 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2095 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1484 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1550 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1566 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1587 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1603 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1609 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1737 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1764 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1776 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1847 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1849 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1862 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1874 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1913 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1998 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2010 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2025 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2037 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1482 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1494 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1506 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1555 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1607 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1611 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1619 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1631 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1650 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1661 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1673 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1717 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1729 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1741 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1773 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1787 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1803 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1814 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1865 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1957 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1969 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1975 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1989 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2001 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2007 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1522 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1530 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1641 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1718 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1770 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1774 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1779 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1791 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1803 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1815 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1823 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1939 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1951 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1959 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1971 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1987 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1999 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2027 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2039 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2051 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_2063 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1577 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1627 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1667 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1677 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1717 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1733 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1837 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1859 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1871 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1913 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1921 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1941 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2054 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2078 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_2090 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_2098 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1520 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1544 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1591 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1608 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1620 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1636 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1662 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1674 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1691 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1716 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1728 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1751 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1829 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1863 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1890 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1902 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1932 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1944 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1956 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1961 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1967 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1971 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1991 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2013 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_2025 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2033 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2048 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1446 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1478 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1502 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1514 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1550 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1556 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1608 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1620 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1638 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1646 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1688 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1891 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1903 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1432 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1443 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1533 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1545 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1602 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1622 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1631 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1671 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1773 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1802 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1873 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1881 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1890 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1929 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1950 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1997 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2005 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2025 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2037 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1483 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1502 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1541 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1606 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1666 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1686 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1720 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1732 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1744 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1756 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1779 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1787 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1796 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1804 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1831 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1855 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1867 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1931 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1499 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1673 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1705 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1847 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1863 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1929 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1935 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1973 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1990 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2002 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2031 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2055 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1338 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1416 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1456 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1556 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1568 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1580 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1592 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1609 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1617 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1629 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1721 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1833 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1839 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1945 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1979 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1989 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2001 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2007 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2145 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1432 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1452 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1477 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1537 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1565 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1582 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1606 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1618 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1647 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1655 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1667 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1693 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1701 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1751 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1774 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1803 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1815 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1827 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1861 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1919 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1943 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1961 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1969 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1981 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2005 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1340 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1439 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1516 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1528 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1532 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1541 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1568 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1580 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1594 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1615 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1658 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1662 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1667 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1684 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1720 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1732 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1740 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1762 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1783 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1799 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1830 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1854 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1866 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1891 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1911 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1524 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1536 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1548 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1581 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1773 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1781 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1799 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1807 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1861 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1929 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1961 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_2011 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1807 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1833 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1839 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1901 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1929 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1951 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1963 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1989 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2001 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2007 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2031 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1524 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1539 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1551 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1593 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1632 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1644 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1654 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1667 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1717 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1721 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1734 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1829 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1837 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1863 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1903 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1920 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1932 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1944 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1984 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1996 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1447 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1459 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1476 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1576 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1614 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1626 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1632 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1636 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1677 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1691 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1723 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1734 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1746 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1765 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1792 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1889 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1901 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1927 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1438 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1549 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1557 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1598 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1606 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1618 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1668 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1686 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1749 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1757 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1764 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1776 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1900 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1913 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1288 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1456 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1476 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1536 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1552 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1576 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1606 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1690 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1720 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1732 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1744 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1783 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1802 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1815 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1819 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1832 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1844 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1860 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1872 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1891 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1915 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1927 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1479 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1523 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1649 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1681 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1708 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1720 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1737 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1764 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1776 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1834 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1863 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1875 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1879 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1929 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1941 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2015 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2027 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2039 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2051 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_2063 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1482 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1512 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1603 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1609 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1615 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1619 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1631 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1635 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1639 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1651 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1661 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1931 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1933 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1939 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1952 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1964 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1989 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2001 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2019 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2035 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1368 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1479 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1681 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1708 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1720 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1732 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1847 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1863 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1903 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1961 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1973 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1979 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1565 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1571 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1609 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1615 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1628 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1640 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1749 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1803 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1815 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1833 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1851 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1891 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1914 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1309 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1526 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1567 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1575 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1579 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1603 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1622 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1634 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1641 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1662 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1674 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1681 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1720 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1732 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1743 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1768 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1830 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1900 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1959 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1990 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2002 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1447 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1517 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1529 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1562 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1574 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1594 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1597 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1605 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1624 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1636 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1765 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1792 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1808 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1835 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1843 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1858 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1870 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1884 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1945 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1971 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_2001 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2028 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_2040 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1284 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1550 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1562 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1584 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1596 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1608 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1620 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1643 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1655 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1660 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1668 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1716 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1805 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1862 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1874 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1886 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1898 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1915 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1935 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1951 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1985 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1552 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1576 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1720 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1763 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1776 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1865 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1877 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1889 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1904 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1920 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1928 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1943 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1955 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1967 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1979 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1365 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1453 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1511 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1581 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1603 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1610 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1622 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1629 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1658 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1761 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1791 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1808 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1820 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1828 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1842 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1849 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1857 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1872 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1884 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1520 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1637 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1659 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1667 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1680 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1692 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1720 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1744 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1779 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1817 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1821 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1827 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1851 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2003 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2027 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1392 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1556 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1587 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1633 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1656 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1929 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1941 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1945 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1958 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1971 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1983 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1996 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_2007 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1528 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1551 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1571 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1577 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1614 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1626 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1638 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1669 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1679 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1687 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1696 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1875 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1904 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1940 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1508 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1873 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1896 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1496 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1508 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1520 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1528 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1677 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1689 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1695 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1734 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1783 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1808 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1831 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1844 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1853 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1870 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1902 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1906 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1960 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1972 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1984 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1412 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1420 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1574 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1586 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1598 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1610 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1620 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1703 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1737 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1764 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1802 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1810 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1823 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1849 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1857 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1878 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1890 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1917 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1929 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1950 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1958 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1961 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1983 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1995 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1446 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1555 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1573 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1604 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1615 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1620 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1636 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1643 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1667 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1679 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1777 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1789 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1957 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1974 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1985 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2007 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2019 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2031 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1332 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1533 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1587 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1639 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1651 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1676 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1706 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1718 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1747 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1759 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1771 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1783 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1847 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1859 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1871 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1883 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1985 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2127 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2135 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_2138 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1498 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1534 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1548 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1584 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1608 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1620 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1644 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1692 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1779 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1783 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1875 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1906 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1918 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1928 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1431 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1602 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1749 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1757 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1789 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1808 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1900 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1919 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1935 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1971 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1983 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1995 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_2007 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1288 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1404 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1521 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1533 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1609 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1631 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1643 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1651 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1677 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1835 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1858 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1901 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1907 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1912 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1933 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1941 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1949 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1953 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1967 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1979 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1531 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1583 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1607 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1648 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1695 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1719 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1829 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1845 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1874 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1886 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1961 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1973 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1979 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1982 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1996 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_2007 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1462 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1482 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1494 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1547 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1573 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1667 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1679 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1683 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1687 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1694 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1706 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1719 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1731 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1743 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1821 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1849 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1866 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1885 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1895 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1907 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2003 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2027 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1510 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1524 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1536 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1542 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1550 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1562 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1581 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1737 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1764 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1776 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1807 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1831 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1873 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1896 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1914 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1938 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1950 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1302 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1614 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1626 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1638 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1673 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1777 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1929 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1942 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1443 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1500 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1543 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1550 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1593 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1612 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1639 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1693 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1701 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1734 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1752 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1760 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1810 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1822 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1832 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1844 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1903 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1911 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1918 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1934 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1942 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1975 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_2011 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1447 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1555 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1587 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1595 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1607 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1619 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1662 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1807 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1819 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1848 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1856 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1895 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1907 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1919 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1928 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1951 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1963 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1325 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1583 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1637 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1735 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1751 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1759 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1847 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1877 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1895 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1403 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1462 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1528 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1550 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1559 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1571 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1579 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1690 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1733 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1828 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1852 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1864 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1885 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1930 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1947 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1971 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1679 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1685 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1689 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1703 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1727 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1735 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1751 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1763 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1771 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1803 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1815 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1827 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1903 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1911 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1918 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1942 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1954 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1971 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1983 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1995 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_2007 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1300 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1444 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1456 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1464 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1565 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1608 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1649 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1658 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1670 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1682 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1777 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1795 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1931 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1942 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1950 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1963 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1979 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1606 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1618 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1644 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1710 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1847 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1867 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1879 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1900 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1905 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1393 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1584 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1639 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1661 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1684 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1696 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1819 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1836 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1847 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1851 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1864 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1897 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1322 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1415 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1527 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1535 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1634 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1646 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1658 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1717 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1721 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1737 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1764 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1849 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1857 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1350 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1550 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1562 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1609 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1667 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1733 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1745 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1492 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1583 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1595 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1744 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1768 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1776 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1793 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1820 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1832 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1844 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1941 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1949 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1689 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1697 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1706 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1787 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1799 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1805 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1830 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1838 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1845 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1857 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1874 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1897 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1907 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1915 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1933 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1500 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1625 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1718 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1730 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1764 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1776 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1829 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1833 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1849 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1863 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1881 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1889 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1902 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1938 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1394 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1406 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1499 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1555 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1579 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1621 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1633 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1694 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1733 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1745 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1749 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1885 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1421 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1432 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1566 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1735 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1746 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1768 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1597 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1616 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1628 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1638 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1675 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1687 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1718 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1754 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1762 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1765 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1773 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1788 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1792 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1831 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1843 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1855 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1867 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1593 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1620 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1639 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1681 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1693 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1699 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1712 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1728 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1757 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1769 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1807 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1811 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1824 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1903 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1923 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1935 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1395 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1495 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1584 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1721 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1725 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1748 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1760 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1860 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1872 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1891 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1903 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1919 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1421 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1471 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1495 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1581 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1587 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1690 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1714 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1776 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1829 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1841 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1863 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1886 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1480 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1504 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1515 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1523 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1555 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1562 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1574 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1649 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1663 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1688 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1721 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1743 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1833 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1845 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1853 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1862 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1874 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1888 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1900 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1912 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1532 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1542 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1550 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1604 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1622 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1643 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1656 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1672 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1687 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1695 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1735 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1743 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1756 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1768 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1793 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1813 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1331 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1386 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1398 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1706 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1752 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1780 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1792 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1808 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1831 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1843 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1855 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1867 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1887 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1907 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1306 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1415 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1432 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1478 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1695 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1805 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1830 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1842 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1863 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1890 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1919 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1943 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1560 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1570 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1580 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1592 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1651 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1662 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1674 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1719 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1725 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1783 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1795 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1807 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1845 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1865 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1873 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1891 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1915 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1927 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1368 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1490 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1510 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1543 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1555 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1590 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1602 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1636 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1660 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1749 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1764 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1772 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1847 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1863 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1387 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1494 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1506 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1538 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1563 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1575 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1588 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1603 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1616 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1628 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1634 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1638 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1669 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1763 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1807 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1819 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1832 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1844 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1856 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1367 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1471 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1596 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1602 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1622 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1650 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1666 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1677 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1699 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1711 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1757 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1793 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1418 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1605 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1627 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1639 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1651 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1657 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1672 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1697 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1713 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1835 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1859 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1871 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1677 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1705 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1717 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1723 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2120 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1704 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1716 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1704 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1716 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_2144 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1680 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1680 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1704 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1716 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1704 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1716 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1704 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1716 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2120 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_2138 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2140 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2128 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2140 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2120 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1691 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1703 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2140 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1764 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1820 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1876 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1908 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1932 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1944 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1988 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2000 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2020 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2032 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2044 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2056 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2088 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2100 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2112 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2132 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1686 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1724 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1736 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1748 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1768 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1824 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1848 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1860 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1904 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1916 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1936 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1960 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1992 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2016 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2048 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2060 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2072 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2128 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_292_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_2129 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_2137 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_296_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_298_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_310_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_314_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_2145 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_320_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_330_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_2125 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_2131 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_2134 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_2138 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_2144 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_2137 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_2145 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_2145 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_2145 ();
endmodule

